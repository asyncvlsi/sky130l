magic
tech sky130l
timestamp 1659178075
<< ndiffusion >>
rect 21 17 26 20
rect 21 14 22 17
rect 25 14 26 17
rect 21 11 26 14
rect 21 8 22 11
rect 25 8 26 11
rect 21 5 26 8
rect 28 5 31 20
rect 33 5 38 20
rect 40 17 45 20
rect 40 14 41 17
rect 44 14 45 17
rect 40 11 45 14
rect 51 16 56 18
rect 51 13 52 16
rect 55 13 56 16
rect 51 12 56 13
rect 58 12 63 18
rect 91 16 96 18
rect 91 13 92 16
rect 95 13 96 16
rect 91 12 96 13
rect 100 16 106 18
rect 100 13 102 16
rect 105 13 106 16
rect 100 12 106 13
rect 40 8 41 11
rect 44 8 45 11
rect 40 5 45 8
<< ndc >>
rect 22 14 25 17
rect 22 8 25 11
rect 41 14 44 17
rect 52 13 55 16
rect 92 13 95 16
rect 102 13 105 16
rect 41 8 44 11
<< ntransistor >>
rect 26 5 28 20
rect 31 5 33 20
rect 38 5 40 20
rect 56 12 58 18
rect 63 12 91 18
rect 96 12 100 18
<< pdiffusion >>
rect 91 35 96 39
rect 51 34 56 35
rect 26 32 31 33
rect 26 29 27 32
rect 30 29 31 32
rect 26 27 31 29
rect 33 32 38 33
rect 33 29 34 32
rect 37 29 38 32
rect 51 31 52 34
rect 55 31 56 34
rect 51 29 56 31
rect 58 29 70 35
rect 84 34 96 35
rect 84 31 86 34
rect 89 31 92 34
rect 95 31 96 34
rect 84 29 96 31
rect 100 34 106 39
rect 100 31 102 34
rect 105 31 106 34
rect 100 29 106 31
rect 33 27 38 29
<< pdc >>
rect 27 29 30 32
rect 34 29 37 32
rect 52 31 55 34
rect 86 31 89 34
rect 92 31 95 34
rect 102 31 105 34
<< ptransistor >>
rect 31 27 33 33
rect 56 29 58 35
rect 70 29 84 35
rect 96 29 100 39
<< polysilicon >>
rect 26 44 37 45
rect 26 41 27 44
rect 30 41 33 44
rect 36 41 37 44
rect 26 40 37 41
rect 70 42 84 43
rect 31 33 33 40
rect 70 39 71 42
rect 74 39 77 42
rect 80 39 84 42
rect 96 39 100 41
rect 56 35 58 37
rect 70 35 84 39
rect 26 20 28 22
rect 31 20 33 27
rect 38 20 40 22
rect 56 18 58 29
rect 70 27 84 29
rect 96 26 100 29
rect 94 25 100 26
rect 94 22 95 25
rect 98 22 100 25
rect 94 21 100 22
rect 63 18 91 20
rect 96 18 100 21
rect 26 0 28 5
rect 31 3 33 5
rect 38 2 40 5
rect 56 2 58 12
rect 63 9 91 12
rect 96 10 100 12
rect 63 6 64 9
rect 67 6 70 9
rect 73 6 76 9
rect 79 6 82 9
rect 85 6 91 9
rect 63 5 91 6
rect 36 1 47 2
rect 21 -1 32 0
rect 21 -4 22 -1
rect 25 -4 28 -1
rect 31 -4 32 -1
rect 36 -2 37 1
rect 40 -2 43 1
rect 46 -2 47 1
rect 36 -3 47 -2
rect 51 1 62 2
rect 51 -2 52 1
rect 55 -2 58 1
rect 61 -2 62 1
rect 51 -3 62 -2
rect 21 -5 32 -4
<< pc >>
rect 27 41 30 44
rect 33 41 36 44
rect 71 39 74 42
rect 77 39 80 42
rect 95 22 98 25
rect 64 6 67 9
rect 70 6 73 9
rect 76 6 79 9
rect 82 6 85 9
rect 22 -4 25 -1
rect 28 -4 31 -1
rect 37 -2 40 1
rect 43 -2 46 1
rect 52 -2 55 1
rect 58 -2 61 1
<< m1 >>
rect 26 41 27 44
rect 30 41 33 44
rect 36 41 37 44
rect 61 39 71 42
rect 74 39 77 42
rect 80 39 81 42
rect 52 34 55 35
rect 27 32 30 33
rect 27 28 30 29
rect 34 32 37 33
rect 34 25 37 29
rect 52 25 55 31
rect 61 31 66 39
rect 102 34 105 35
rect 85 31 86 34
rect 89 31 92 34
rect 95 31 96 34
rect 61 28 62 31
rect 65 28 66 31
rect 34 22 95 25
rect 98 22 99 25
rect 22 17 25 18
rect 22 11 25 14
rect 22 7 25 8
rect 41 17 44 22
rect 41 11 44 14
rect 52 16 55 22
rect 52 12 55 13
rect 78 16 79 19
rect 82 16 85 19
rect 88 16 89 19
rect 92 16 95 17
rect 78 9 86 16
rect 92 12 95 13
rect 102 16 105 31
rect 41 7 44 8
rect 63 6 64 9
rect 67 6 70 9
rect 73 6 76 9
rect 79 6 82 9
rect 85 6 86 9
rect 102 1 105 13
rect 21 -4 22 -1
rect 25 -4 28 -1
rect 31 -4 32 -1
rect 36 -2 37 1
rect 40 -2 43 1
rect 46 -2 47 1
rect 51 -2 52 1
rect 55 -2 58 1
rect 61 -2 105 1
<< m2c >>
rect 62 28 65 31
rect 79 16 82 19
rect 85 16 88 19
<< m2 >>
rect 26 34 96 37
rect 26 28 31 34
rect 61 31 66 32
rect 61 28 62 31
rect 65 28 66 31
rect 21 13 26 18
rect 61 13 66 28
rect 78 30 96 34
rect 78 19 89 30
rect 78 16 79 19
rect 82 16 85 19
rect 88 16 89 19
rect 78 15 89 16
rect 91 13 96 17
rect 21 10 96 13
rect 21 7 26 10
<< labels >>
rlabel ndiffusion 25 6 25 6 7 GND
rlabel polysilicon 27 21 27 21 7 in(0)
rlabel pdiffusion 30 28 30 28 7 Vdd
rlabel polysilicon 32 21 32 21 7 in(1)
rlabel polysilicon 32 26 32 26 7 in(1)
rlabel pdiffusion 37 28 37 28 7 out
rlabel polysilicon 39 21 39 21 7 in(2)
rlabel ndiffusion 44 6 44 6 7 out
rlabel ndiffusion 102 13 102 13 3 #10
rlabel pdiffusion 105 30 105 30 7 #10
rlabel polysilicon 97 19 97 19 3 out
rlabel ndiffusion 92 13 92 13 3 GND
rlabel polysilicon 64 19 64 19 3 Vdd
rlabel ndiffusion 59 13 59 13 3 #12
rlabel polysilicon 57 19 57 19 3 #10
rlabel ndiffusion 52 13 52 13 3 out
rlabel polysilicon 83 28 83 28 7 GND
rlabel pdiffusion 69 30 69 30 7 #11
rlabel pdiffusion 62 30 62 30 7 out
rlabel polysilicon 57 28 57 28 7 #10
rlabel pdiffusion 55 30 55 30 7 #11
rlabel polysilicon 99 28 99 28 7 out
rlabel pdiffusion 95 30 95 30 7 Vdd
flabel m2 26 34 96 37 0 FreeSans 11 0 0 0 Vdd
port 1 nsew
flabel m2 22 10 96 13 0 FreeSans 11 0 0 0 GND
flabel m1 21 -4 32 -1 0 FreeSans 11 0 0 0 in(0)
port 3 nsew
flabel m1 26 41 37 44 0 FreeSans 11 0 0 0 in(1)
port 4 nsew
flabel m1 36 -2 47 1 0 FreeSans 11 0 0 0 in(2)
port 5 nsew
flabel m1 34 22 99 25 0 FreeSans 11 0 0 0 out
port 6 nsew
<< end >>
