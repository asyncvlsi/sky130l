magic
tech sky130l
timestamp 1639029389
<< ndiffusion >>
rect 8 10 13 16
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 6 20 16
rect 22 15 27 16
rect 22 12 23 15
rect 26 12 27 15
rect 22 6 27 12
rect 34 15 39 16
rect 34 12 35 15
rect 38 12 39 15
rect 34 10 39 12
rect 41 14 48 16
rect 41 11 43 14
rect 46 11 48 14
rect 41 10 48 11
rect 44 6 48 10
rect 50 10 55 16
rect 50 7 51 10
rect 54 7 55 10
rect 50 6 55 7
rect 62 15 67 16
rect 62 12 63 15
rect 66 12 67 15
rect 62 6 67 12
rect 69 10 74 16
rect 69 7 70 10
rect 73 7 74 10
rect 69 6 74 7
<< ndc >>
rect 9 7 12 10
rect 23 12 26 15
rect 35 12 38 15
rect 43 11 46 14
rect 51 7 54 10
rect 63 12 66 15
rect 70 7 73 10
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
rect 39 10 41 16
rect 48 6 50 16
rect 67 6 69 16
<< pdiffusion >>
rect 8 37 13 38
rect 8 34 9 37
rect 12 34 13 37
rect 8 23 13 34
rect 15 31 19 38
rect 15 30 20 31
rect 15 27 16 30
rect 19 27 20 30
rect 15 23 20 27
rect 22 27 27 31
rect 22 24 23 27
rect 26 24 27 27
rect 22 23 27 24
rect 34 27 39 38
rect 34 24 35 27
rect 38 24 39 27
rect 34 23 39 24
rect 41 23 48 38
rect 50 33 55 38
rect 50 30 51 33
rect 54 30 55 33
rect 50 23 55 30
rect 62 37 67 38
rect 62 34 63 37
rect 66 34 67 37
rect 62 23 67 34
rect 69 27 74 38
rect 69 24 70 27
rect 73 24 74 27
rect 69 23 74 24
<< pdc >>
rect 9 34 12 37
rect 16 27 19 30
rect 23 24 26 27
rect 35 24 38 27
rect 51 30 54 33
rect 63 34 66 37
rect 70 24 73 27
<< ptransistor >>
rect 13 23 15 38
rect 20 23 22 31
rect 39 23 41 38
rect 48 23 50 38
rect 67 23 69 38
<< polysilicon >>
rect 10 45 15 46
rect 10 42 11 45
rect 14 42 15 45
rect 10 41 15 42
rect 13 38 15 41
rect 20 45 25 46
rect 20 42 21 45
rect 24 42 25 45
rect 20 41 25 42
rect 36 45 41 46
rect 36 42 37 45
rect 40 42 41 45
rect 36 41 41 42
rect 20 31 22 41
rect 39 38 41 41
rect 48 45 53 46
rect 48 42 49 45
rect 52 42 53 45
rect 48 41 53 42
rect 67 45 72 46
rect 67 42 68 45
rect 71 42 72 45
rect 67 41 72 42
rect 48 38 50 41
rect 67 38 69 41
rect 13 16 15 23
rect 20 16 22 23
rect 39 16 41 23
rect 48 16 50 23
rect 67 16 69 23
rect 39 8 41 10
rect 13 4 15 6
rect 20 4 22 6
rect 48 4 50 6
rect 67 4 69 6
<< pc >>
rect 11 42 14 45
rect 21 42 24 45
rect 37 42 40 45
rect 49 42 52 45
rect 68 42 71 45
<< m1 >>
rect 10 45 15 46
rect 10 42 11 45
rect 14 42 15 45
rect 20 45 41 46
rect 20 42 21 45
rect 24 42 37 45
rect 40 42 41 45
rect 48 45 53 46
rect 48 42 49 45
rect 52 42 53 45
rect 62 45 72 46
rect 62 42 63 45
rect 66 42 68 45
rect 71 42 72 45
rect 9 37 66 39
rect 8 34 9 37
rect 12 36 63 37
rect 12 34 13 36
rect 63 33 66 34
rect 16 30 51 33
rect 54 30 55 33
rect 70 27 73 28
rect 16 26 19 27
rect 22 24 23 27
rect 26 24 27 27
rect 34 24 35 27
rect 38 24 39 27
rect 35 21 38 24
rect 70 21 73 24
rect 23 19 73 21
rect 26 18 73 19
rect 23 15 26 16
rect 63 15 66 18
rect 22 12 23 15
rect 26 12 27 15
rect 34 12 35 15
rect 38 12 39 15
rect 43 14 46 15
rect 62 12 63 15
rect 66 12 67 15
rect 8 7 9 10
rect 12 9 13 10
rect 43 9 46 11
rect 70 10 74 11
rect 12 7 46 9
rect 8 6 46 7
rect 50 7 51 10
rect 54 9 55 10
rect 54 7 70 9
rect 73 7 74 10
rect 50 6 74 7
rect 22 0 23 3
rect 22 -1 26 0
<< m2c >>
rect 63 42 66 45
rect 27 24 30 27
rect 23 16 26 19
rect 31 12 34 15
rect 23 0 26 3
<< m2 >>
rect 62 45 67 46
rect 62 43 63 45
rect 30 42 63 43
rect 66 42 67 45
rect 30 41 67 42
rect 30 28 32 41
rect 26 27 32 28
rect 26 24 27 27
rect 30 24 32 27
rect 26 23 32 24
rect 22 19 27 20
rect 22 16 23 19
rect 26 16 27 19
rect 22 15 27 16
rect 25 4 27 15
rect 30 16 32 23
rect 30 15 35 16
rect 30 12 31 15
rect 34 12 35 15
rect 30 11 35 12
rect 22 3 27 4
rect 22 0 23 3
rect 26 0 27 3
rect 22 -1 27 0
<< labels >>
rlabel ndiffusion 23 7 23 7 3 Y
rlabel polysilicon 14 17 14 17 3 A
rlabel polysilicon 14 22 14 22 3 A
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 24 9 24 3 #5
rlabel ndiffusion 51 7 51 7 3 #10
rlabel polysilicon 49 17 49 17 3 B
rlabel polysilicon 49 22 49 22 3 B
rlabel ndiffusion 42 11 42 11 3 GND
rlabel pdiffusion 35 24 35 24 3 Y
rlabel ndiffusion 70 7 70 7 3 #10
rlabel pdiffusion 70 24 70 24 3 Y
rlabel ndiffusion 63 7 63 7 3 Y
rlabel pdiffusion 63 24 63 24 3 #5
rlabel pdiffusion 16 24 16 24 3 Vdd
rlabel pdiffusion 51 24 51 24 3 Vdd
rlabel m1 11 43 11 43 3 A
port 6 e
rlabel m1 49 43 49 43 3 B
port 4 e
rlabel m1 27 31 27 31 3 Vdd
port 2 e
rlabel m1 31 7 31 7 3 GND
port 1 e
rlabel m1 23 0 23 0 3 Y
port 5 e
rlabel polysilicon 68 17 68 17 3 _S
rlabel polysilicon 68 22 68 22 3 _S
rlabel polysilicon 21 17 21 17 3 S
rlabel polysilicon 21 22 21 22 3 S
rlabel polysilicon 40 17 40 17 3 S
rlabel polysilicon 40 22 40 22 3 S
rlabel pc 38 43 38 43 3 S
port 3 e
rlabel pdiffusion 23 24 23 24 3 _S
rlabel ndiffusion 35 11 35 11 3 _S
<< end >>
