magic
tech sky130l
timestamp 1635619534
<< ndiffusion >>
rect 6 10 11 12
rect 6 7 7 10
rect 10 7 11 10
rect 6 4 11 7
rect 13 11 20 12
rect 13 8 15 11
rect 18 8 20 11
rect 13 4 20 8
rect 22 10 27 12
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
rect 29 11 34 12
rect 29 8 30 11
rect 33 8 34 11
rect 29 6 34 8
rect 22 4 26 6
<< ndc >>
rect 7 7 10 10
rect 15 8 18 11
rect 23 7 26 10
rect 30 8 33 11
<< ntransistor >>
rect 11 4 13 12
rect 20 4 22 12
rect 27 6 29 12
<< pdiffusion >>
rect 6 23 11 25
rect 6 20 7 23
rect 10 20 11 23
rect 6 19 11 20
rect 15 23 20 25
rect 15 20 16 23
rect 19 20 20 23
rect 15 19 20 20
rect 24 23 29 25
rect 24 20 25 23
rect 28 20 29 23
rect 24 19 29 20
<< pdc >>
rect 7 20 10 23
rect 16 20 19 23
rect 25 20 28 23
<< ptransistor >>
rect 11 19 15 25
rect 20 19 24 25
<< polysilicon >>
rect 10 32 15 33
rect 10 29 11 32
rect 14 29 15 32
rect 10 28 15 29
rect 11 25 15 28
rect 20 25 24 27
rect 11 17 15 19
rect 20 17 24 19
rect 11 12 13 17
rect 20 12 22 17
rect 27 12 29 14
rect 11 2 13 4
rect 20 2 22 4
rect 27 2 29 6
rect 19 1 24 2
rect 19 -2 20 1
rect 23 -2 24 1
rect 19 -3 24 -2
rect 27 1 32 2
rect 27 -2 28 1
rect 31 -2 32 1
rect 27 -3 32 -2
<< pc >>
rect 11 29 14 32
rect 20 -2 23 1
rect 28 -2 31 1
<< m1 >>
rect 10 29 11 32
rect 14 29 27 32
rect 7 23 10 24
rect 7 10 10 20
rect 16 23 19 25
rect 24 24 27 29
rect 16 19 19 20
rect 23 23 29 24
rect 23 20 25 23
rect 28 20 29 23
rect 23 19 29 20
rect 15 11 18 12
rect 15 7 18 8
rect 23 10 26 19
rect 7 1 10 7
rect 23 6 26 7
rect 30 11 33 12
rect 30 6 33 8
rect 7 -2 20 1
rect 23 -2 24 1
rect 27 -2 28 1
rect 31 -2 32 1
<< m2c >>
rect 16 20 19 23
rect 15 8 18 11
rect 30 8 33 11
<< m2 >>
rect 11 23 22 24
rect 11 20 16 23
rect 19 20 22 23
rect 11 19 22 20
rect 14 11 34 12
rect 14 8 15 11
rect 18 8 30 11
rect 33 8 34 11
rect 14 7 19 8
rect 29 7 34 8
<< labels >>
rlabel polysilicon 28 13 28 13 3 Reset
rlabel polysilicon 21 13 21 13 3 df
rlabel polysilicon 21 18 21 18 3 df
rlabel polysilicon 12 13 12 13 3 dt
rlabel polysilicon 12 18 12 18 3 dt
rlabel pdc 9 21 9 21 3 df
rlabel ndc 8 9 8 9 3 df
rlabel ndc 24 9 24 9 3 dt
rlabel ndc 16 9 16 9 3 GND
rlabel pdc 26 21 26 21 3 dt
rlabel m1 8 16 8 16 3 df
rlabel m1 24 15 24 15 1 dt
rlabel m2c 31 9 31 9 7 GND
rlabel m1 17 24 17 24 1 Vdd
rlabel m2 13 21 13 21 1 Vdd
<< end >>
