magic
tech sky130l
timestamp 1639252531
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 11 20 12
rect 15 8 16 11
rect 19 8 20 11
rect 15 6 20 8
rect 22 10 27 12
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
rect 29 11 34 12
rect 29 8 30 11
rect 33 8 34 11
rect 29 6 34 8
<< ndc >>
rect 9 7 12 10
rect 16 8 19 11
rect 23 7 26 10
rect 30 8 33 11
<< ntransistor >>
rect 13 6 15 12
rect 20 6 22 12
rect 27 6 29 12
<< pdiffusion >>
rect 8 37 13 42
rect 8 34 9 37
rect 12 34 13 37
rect 8 19 13 34
rect 15 19 20 42
rect 22 19 27 42
rect 29 23 34 42
rect 29 20 30 23
rect 33 20 34 23
rect 29 19 34 20
<< pdc >>
rect 9 34 12 37
rect 30 20 33 23
<< ptransistor >>
rect 13 19 15 42
rect 20 19 22 42
rect 27 19 29 42
<< polysilicon >>
rect 10 49 15 50
rect 10 46 11 49
rect 14 46 15 49
rect 10 45 15 46
rect 18 49 23 50
rect 18 46 19 49
rect 22 46 23 49
rect 18 45 23 46
rect 26 49 31 50
rect 26 46 27 49
rect 30 46 31 49
rect 26 45 31 46
rect 13 42 15 45
rect 20 42 22 45
rect 27 42 29 45
rect 13 12 15 19
rect 20 12 22 19
rect 27 12 29 19
rect 13 4 15 6
rect 20 4 22 6
rect 27 4 29 6
<< pc >>
rect 11 46 14 49
rect 19 46 22 49
rect 27 46 30 49
<< m1 >>
rect 11 49 15 50
rect 14 46 15 49
rect 11 45 15 46
rect 19 49 23 50
rect 22 46 23 49
rect 19 45 23 46
rect 27 49 31 50
rect 30 46 31 49
rect 27 45 31 46
rect 9 37 12 38
rect 9 33 12 34
rect 30 23 33 24
rect 15 12 18 20
rect 15 11 19 12
rect 30 11 33 20
rect 9 10 12 11
rect 15 8 16 11
rect 15 7 19 8
rect 23 10 27 11
rect 26 7 27 10
rect 9 6 12 7
rect 23 6 27 7
rect 30 6 33 8
<< m2c >>
rect 9 34 12 37
rect 15 20 18 23
rect 30 20 33 23
rect 9 7 12 10
rect 23 7 26 10
<< m2 >>
rect 8 37 33 38
rect 8 34 9 37
rect 12 34 33 37
rect 8 33 33 34
rect 14 23 34 24
rect 14 20 15 23
rect 18 22 30 23
rect 18 20 19 22
rect 14 19 19 20
rect 29 20 30 22
rect 33 20 34 23
rect 29 19 34 20
rect 8 10 27 11
rect 8 7 9 10
rect 12 7 23 10
rect 26 7 27 10
rect 8 6 27 7
<< labels >>
rlabel ndiffusion 30 7 30 7 3 Y
rlabel pdiffusion 30 20 30 20 3 Y
rlabel polysilicon 28 13 28 13 3 C
rlabel polysilicon 28 18 28 18 3 C
rlabel ndiffusion 23 7 23 7 3 GND
rlabel polysilicon 21 13 21 13 3 B
rlabel polysilicon 21 18 21 18 3 B
rlabel ndiffusion 16 7 16 7 3 Y
rlabel polysilicon 14 13 14 13 3 A
rlabel polysilicon 14 18 14 18 3 A
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 20 9 20 3 Vdd
rlabel pc 12 47 12 47 3 A
port 6 e
rlabel pc 20 47 20 47 3 B
port 4 e
rlabel pc 28 47 28 47 3 C
port 3 e
rlabel m1 10 34 10 34 3 Vdd
port 2 e
rlabel m2c 17 21 17 21 1 Y
rlabel ndc 10 8 10 8 3 GND
port 1 e
<< end >>
