magic
tech sky130l
timestamp 1639177113
<< ndiffusion >>
rect 8 10 13 16
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 6 20 16
rect 22 15 27 16
rect 22 12 23 15
rect 26 12 27 15
rect 22 6 27 12
<< ndc >>
rect 9 7 12 10
rect 23 12 26 15
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
<< pdiffusion >>
rect 8 30 13 31
rect 8 27 9 30
rect 12 27 13 30
rect 8 23 13 27
rect 15 27 20 31
rect 15 24 16 27
rect 19 24 20 27
rect 15 23 20 24
rect 22 30 27 31
rect 22 27 23 30
rect 26 27 27 30
rect 22 23 27 27
<< pdc >>
rect 9 27 12 30
rect 16 24 19 27
rect 23 27 26 30
<< ptransistor >>
rect 13 23 15 31
rect 20 23 22 31
<< polysilicon >>
rect 10 40 15 41
rect 10 37 11 40
rect 14 37 15 40
rect 10 36 15 37
rect 13 31 15 36
rect 20 40 25 41
rect 20 37 21 40
rect 24 37 25 40
rect 20 36 25 37
rect 20 31 22 36
rect 13 16 15 23
rect 20 16 22 23
rect 13 4 15 6
rect 20 4 22 6
<< pc >>
rect 11 37 14 40
rect 21 37 24 40
<< m1 >>
rect 10 40 15 41
rect 10 37 11 40
rect 14 37 15 40
rect 20 40 25 41
rect 20 37 21 40
rect 24 37 25 40
rect 9 30 12 31
rect 5 27 9 30
rect 23 30 27 31
rect 5 26 12 27
rect 15 27 19 28
rect 15 24 16 27
rect 26 27 27 30
rect 23 26 27 27
rect 15 23 19 24
rect 15 17 18 23
rect 23 15 26 16
rect 9 10 12 11
rect 9 6 12 7
rect 23 1 26 12
<< m2c >>
rect 9 27 12 30
rect 23 27 26 30
rect 15 14 18 17
rect 23 12 26 15
rect 9 7 12 10
<< m2 >>
rect 8 30 13 31
rect 8 27 9 30
rect 12 28 13 30
rect 22 30 27 31
rect 22 28 23 30
rect 12 27 23 28
rect 26 27 27 30
rect 8 26 27 27
rect 14 17 27 18
rect 14 14 15 17
rect 18 16 27 17
rect 18 14 19 16
rect 14 13 19 14
rect 22 15 27 16
rect 22 12 23 15
rect 26 12 27 15
rect 22 11 27 12
rect 8 10 13 11
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
<< labels >>
rlabel ndiffusion 23 7 23 7 3 Y
rlabel pdiffusion 23 24 23 24 3 Vdd
rlabel polysilicon 21 17 21 17 3 B
rlabel polysilicon 21 22 21 22 3 B
rlabel pdiffusion 16 24 16 24 3 Y
rlabel polysilicon 14 22 14 22 3 A
rlabel pdiffusion 9 24 9 24 3 Vdd
rlabel m1 21 38 21 38 3 B
port 3 e
rlabel m1 11 38 11 38 3 A
port 5 e
rlabel m1 6 27 6 27 3 Vdd
port 2 e
rlabel m1 24 2 24 2 3 Y
port 4 e
rlabel m1 10 7 10 7 3 GND
port 1 e
rlabel polysilicon 14 17 14 17 3 A
<< end >>
