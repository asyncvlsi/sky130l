magic
tech sky130l
timestamp 1636659416
<< ndiffusion >>
rect 7 11 12 12
rect 7 8 8 11
rect 11 8 12 11
rect 7 6 12 8
rect 14 6 19 12
rect 21 11 26 12
rect 21 8 22 11
rect 25 8 26 11
rect 21 6 26 8
<< ndc >>
rect 8 8 11 11
rect 22 8 25 11
<< ntransistor >>
rect 12 6 14 12
rect 19 6 21 12
<< pdiffusion >>
rect 7 23 12 31
rect 7 20 8 23
rect 11 20 12 23
rect 7 19 12 20
rect 14 19 19 31
rect 21 23 26 31
rect 21 20 22 23
rect 25 20 26 23
rect 21 19 26 20
<< pdc >>
rect 8 20 11 23
rect 22 20 25 23
<< ptransistor >>
rect 12 19 14 31
rect 19 19 21 31
<< polysilicon >>
rect 12 31 14 33
rect 19 31 21 33
rect 12 12 14 19
rect 19 12 21 19
rect 12 4 14 6
rect 7 3 14 4
rect 7 0 8 3
rect 11 2 14 3
rect 19 4 21 6
rect 19 3 26 4
rect 19 2 22 3
rect 11 0 12 2
rect 7 -1 12 0
rect 21 0 22 2
rect 25 0 26 3
rect 21 -1 26 0
<< pc >>
rect 8 0 11 3
rect 22 0 25 3
<< m1 >>
rect 8 23 11 24
rect 22 23 25 24
rect 8 19 11 20
rect 8 11 11 12
rect 8 7 11 8
rect 7 3 12 4
rect 7 0 8 3
rect 11 0 12 3
rect 7 -1 12 0
rect 9 -4 12 -1
rect 15 -4 18 20
rect 22 19 25 20
rect 22 11 25 12
rect 22 7 25 8
rect 21 3 26 4
rect 21 0 22 3
rect 25 0 26 3
rect 21 -1 26 0
rect 21 -4 24 -1
<< m2c >>
rect 8 20 11 23
rect 15 20 18 23
rect 8 8 11 11
rect 22 20 25 23
rect 22 8 25 11
<< m2 >>
rect 7 23 12 24
rect 7 20 8 23
rect 11 20 12 23
rect 0 18 12 20
rect 14 23 26 24
rect 14 20 15 23
rect 18 22 22 23
rect 18 20 19 22
rect 14 19 19 20
rect 21 20 22 22
rect 25 20 26 23
rect 21 19 26 20
rect 21 12 33 14
rect 7 11 26 12
rect 7 8 8 11
rect 11 10 22 11
rect 11 8 12 10
rect 7 7 12 8
rect 21 8 22 10
rect 25 8 26 11
rect 21 7 26 8
<< labels >>
rlabel ndiffusion 22 7 22 7 3 GND
rlabel polysilicon 20 13 20 13 3 in(1)
rlabel polysilicon 20 18 20 18 3 in(1)
rlabel ndiffusion 15 7 15 7 3 out
rlabel polysilicon 13 13 13 13 3 in(0)
rlabel polysilicon 13 18 13 18 3 in(0)
rlabel ndiffusion 8 7 8 7 3 GND
rlabel pdiffusion 8 20 8 20 3 Vdd
rlabel m1 16 1 16 1 3 out
port 4 e
rlabel pdiffusion 22 20 22 20 3 out
rlabel m2 24 13 24 13 3 GND
port 1 e
rlabel m1 10 -2 10 -2 3 in(0)
port 5 e
rlabel m1 23 -2 23 -2 3 in(1)
port 3 e
rlabel m2 0 18 2 20 3 Vdd
rlabel m2 31 12 33 14 7 GND
<< end >>
