magic
tech sky130l
timestamp 1636603609
<< ndiffusion >>
rect 8 15 13 16
rect 8 12 9 15
rect 12 12 13 15
rect 8 6 13 12
rect 15 11 20 16
rect 15 8 16 11
rect 19 8 20 11
rect 15 6 20 8
rect 22 6 27 16
rect 29 11 34 16
rect 29 8 30 11
rect 33 8 34 11
rect 29 6 34 8
rect 36 15 41 16
rect 36 12 37 15
rect 40 12 41 15
rect 36 6 41 12
<< ndc >>
rect 9 12 12 15
rect 16 8 19 11
rect 30 8 33 11
rect 37 12 40 15
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
rect 27 6 29 16
rect 34 6 36 16
<< pdiffusion >>
rect 8 33 13 38
rect 8 30 9 33
rect 12 30 13 33
rect 8 23 13 30
rect 15 28 20 38
rect 15 25 16 28
rect 19 25 20 28
rect 15 23 20 25
rect 22 28 27 38
rect 22 25 23 28
rect 26 25 27 28
rect 22 23 27 25
rect 29 28 34 38
rect 29 25 30 28
rect 33 25 34 28
rect 29 23 34 25
rect 36 33 41 38
rect 36 30 37 33
rect 40 30 41 33
rect 36 23 41 30
<< pdc >>
rect 9 30 12 33
rect 16 25 19 28
rect 23 25 26 28
rect 30 25 33 28
rect 37 30 40 33
<< ptransistor >>
rect 13 23 15 38
rect 20 23 22 38
rect 27 23 29 38
rect 34 23 36 38
<< polysilicon >>
rect 10 45 15 46
rect 10 42 11 45
rect 14 42 15 45
rect 10 41 15 42
rect 18 45 23 46
rect 18 42 19 45
rect 22 42 23 45
rect 18 41 23 42
rect 26 45 31 46
rect 26 42 27 45
rect 30 42 31 45
rect 26 41 31 42
rect 34 45 39 46
rect 34 42 35 45
rect 38 42 39 45
rect 34 41 39 42
rect 13 38 15 41
rect 20 38 22 41
rect 27 38 29 41
rect 34 38 36 41
rect 13 16 15 23
rect 20 16 22 23
rect 27 16 29 23
rect 34 16 36 23
rect 13 4 15 6
rect 20 4 22 6
rect 27 4 29 6
rect 34 4 36 6
<< pc >>
rect 11 42 14 45
rect 19 42 22 45
rect 27 42 30 45
rect 35 42 38 45
<< m1 >>
rect 12 46 15 48
rect 10 45 15 46
rect 10 42 11 45
rect 14 42 15 45
rect 10 41 15 42
rect 18 46 21 48
rect 27 46 30 48
rect 36 46 39 48
rect 18 45 23 46
rect 18 42 19 45
rect 22 42 23 45
rect 18 41 23 42
rect 26 45 31 46
rect 26 42 27 45
rect 30 42 31 45
rect 26 41 31 42
rect 34 45 39 46
rect 34 42 35 45
rect 38 42 39 45
rect 34 41 39 42
rect 36 34 39 36
rect 9 33 12 34
rect 9 29 12 30
rect 36 33 40 34
rect 36 30 37 33
rect 36 29 40 30
rect 16 28 19 29
rect 16 24 19 25
rect 23 28 27 29
rect 26 25 27 28
rect 23 24 27 25
rect 30 28 33 29
rect 30 24 33 25
rect 9 15 12 16
rect 24 12 27 24
rect 37 15 40 16
rect 9 11 12 12
rect 15 11 19 12
rect 15 8 16 11
rect 15 7 19 8
rect 22 11 27 12
rect 22 8 23 11
rect 26 8 27 11
rect 22 7 27 8
rect 30 11 33 12
rect 37 11 40 12
rect 15 -14 18 7
rect 30 -1 33 8
rect 32 -4 33 -1
rect 30 -6 33 -4
<< m2c >>
rect 9 30 12 33
rect 37 30 40 33
rect 16 25 19 28
rect 30 25 33 28
rect 9 12 12 15
rect 37 12 40 15
rect 16 8 19 11
rect 23 8 26 11
rect 30 8 33 11
rect 29 -4 32 -1
<< m2 >>
rect -3 33 57 34
rect -3 32 9 33
rect 8 30 9 32
rect 12 32 37 33
rect 12 30 13 32
rect 8 29 13 30
rect 36 30 37 32
rect 40 32 57 33
rect 40 30 41 32
rect 36 29 41 30
rect 15 28 20 29
rect 29 28 34 29
rect 15 25 16 28
rect 19 26 30 28
rect 19 25 20 26
rect 15 24 20 25
rect 29 25 30 26
rect 33 25 34 28
rect 29 24 34 25
rect 8 15 41 16
rect 8 12 9 15
rect 12 14 37 15
rect 12 12 13 14
rect 36 12 37 14
rect 40 12 41 15
rect 8 11 13 12
rect 15 11 20 12
rect 15 8 16 11
rect 19 10 20 11
rect 22 11 27 12
rect 22 10 23 11
rect 19 8 23 10
rect 26 8 27 11
rect 15 7 20 8
rect 22 7 27 8
rect 29 11 34 12
rect 36 11 41 12
rect 29 8 30 11
rect 33 8 34 11
rect 29 7 34 8
rect 27 -1 33 0
rect 27 -4 29 -1
rect 32 -2 33 -1
rect 32 -4 42 -2
rect 27 -6 33 -4
<< labels >>
rlabel ndiffusion 37 7 37 7 3 #3
rlabel polysilicon 35 17 35 17 3 A
rlabel polysilicon 35 22 35 22 3 A
rlabel polysilicon 28 17 28 17 3 C
rlabel polysilicon 28 22 28 22 3 C
rlabel pdiffusion 23 24 23 24 3 Y
rlabel polysilicon 21 17 21 17 3 D
rlabel polysilicon 21 22 21 22 3 D
rlabel polysilicon 14 17 14 17 3 B
rlabel polysilicon 14 22 14 22 3 B
rlabel m1 13 47 13 47 3 B
port 5 e
rlabel m1 28 47 28 47 3 C
port 4 e
rlabel m1 19 47 19 47 3 D
port 3 e
rlabel m1 37 47 37 47 3 A
port 7 e
rlabel pdiffusion 37 35 37 35 3 Vdd
port 2 e
rlabel m1 16 5 16 5 3 Y
port 6 e
rlabel m1 31 5 31 5 3 GND
port 1 e
rlabel pdiffusion 9 30 9 30 3 Vdd
rlabel pdiffusion 17 25 17 25 3 #9
rlabel m2c 31 26 31 26 3 #9
rlabel m2c 31 9 31 9 3 GND
rlabel m2c 17 9 17 9 3 Y
rlabel m2c 10 13 10 13 3 #3
rlabel m2c 38 32 38 32 3 Vdd
<< end >>
