magic
tech sky130l
timestamp 1636154993
<< ndiffusion >>
rect 8 11 13 12
rect 8 8 9 11
rect 12 8 13 11
rect 8 6 13 8
rect 15 11 20 12
rect 15 8 16 11
rect 19 8 20 11
rect 15 6 20 8
rect 22 11 27 12
rect 22 8 23 11
rect 26 8 27 11
rect 22 6 27 8
<< ndc >>
rect 9 8 12 11
rect 16 8 19 11
rect 23 8 26 11
<< ntransistor >>
rect 13 6 15 12
rect 20 6 22 12
<< pdiffusion >>
rect 8 33 13 34
rect 8 30 9 33
rect 12 30 13 33
rect 8 19 13 30
rect 15 19 20 34
rect 22 23 27 34
rect 22 20 23 23
rect 26 20 27 23
rect 22 19 27 20
<< pdc >>
rect 9 30 12 33
rect 23 20 26 23
<< ptransistor >>
rect 13 19 15 34
rect 20 19 22 34
<< polysilicon >>
rect 13 34 15 36
rect 20 34 22 36
rect 13 12 15 19
rect 20 12 22 19
rect 13 3 15 6
rect 20 3 22 6
rect 11 2 16 3
rect 11 -1 12 2
rect 15 -1 16 2
rect 11 -2 16 -1
rect 19 2 24 3
rect 19 -1 20 2
rect 23 -1 24 2
rect 19 -2 24 -1
<< pc >>
rect 12 -1 15 2
rect 20 -1 23 2
<< m1 >>
rect 9 33 12 34
rect 9 29 12 30
rect 23 23 26 24
rect 15 12 18 20
rect 23 19 26 20
rect 9 11 12 12
rect 9 7 12 8
rect 15 11 19 12
rect 15 8 16 11
rect 15 7 19 8
rect 23 11 26 12
rect 23 7 26 8
rect 12 2 15 3
rect 12 -2 15 -1
rect 20 2 24 3
rect 23 -1 24 2
rect 20 -2 24 -1
<< m2c >>
rect 9 30 12 33
rect 15 20 18 23
rect 23 20 26 23
rect 9 8 12 11
rect 23 8 26 11
rect 12 -1 15 2
rect 20 -1 23 2
<< m2 >>
rect 8 33 13 34
rect 8 32 9 33
rect 6 30 9 32
rect 12 30 13 33
rect 8 29 13 30
rect 14 23 19 24
rect 14 20 15 23
rect 18 22 19 23
rect 22 23 27 24
rect 22 22 23 23
rect 18 20 23 22
rect 26 22 27 23
rect 26 20 30 22
rect 14 19 19 20
rect 22 19 27 20
rect 8 11 13 12
rect 8 10 9 11
rect 6 8 9 10
rect 12 10 13 11
rect 22 11 27 12
rect 22 10 23 11
rect 12 8 23 10
rect 26 8 27 11
rect 8 7 13 8
rect 22 7 27 8
rect 11 2 16 3
rect 6 0 12 2
rect 11 -1 12 0
rect 15 -1 16 2
rect 11 -2 16 -1
rect 19 2 24 3
rect 19 -1 20 2
rect 23 0 27 2
rect 23 -1 24 0
rect 19 -2 24 -1
<< labels >>
rlabel m2 7 9 7 9 3 GND
rlabel m2 26 1 26 1 8 B
rlabel m2 8 1 8 1 2 A
rlabel m2 7 31 7 31 4 Vdd
rlabel m2 29 21 29 21 7 Y
<< end >>
