magic
tech sky130l
timestamp 1636172055
<< ndiffusion >>
rect 8 10 13 16
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 15 20 16
rect 15 12 16 15
rect 19 12 20 15
rect 15 6 20 12
rect 22 10 27 16
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
rect 29 10 34 16
rect 29 7 30 10
rect 33 7 34 10
rect 29 6 34 7
rect 36 10 41 16
rect 36 7 37 10
rect 40 7 41 10
rect 36 6 41 7
<< ndc >>
rect 9 7 12 10
rect 16 12 19 15
rect 23 7 26 10
rect 30 7 33 10
rect 37 7 40 10
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
rect 27 6 29 16
rect 34 6 36 16
<< pdiffusion >>
rect 8 28 13 38
rect 8 25 9 28
rect 12 25 13 28
rect 8 23 13 25
rect 15 23 20 38
rect 22 27 27 38
rect 22 24 23 27
rect 26 24 27 27
rect 22 23 27 24
rect 29 23 34 38
rect 36 28 41 38
rect 36 25 37 28
rect 40 25 41 28
rect 36 23 41 25
<< pdc >>
rect 9 25 12 28
rect 23 24 26 27
rect 37 25 40 28
<< ptransistor >>
rect 13 23 15 38
rect 20 23 22 38
rect 27 23 29 38
rect 34 23 36 38
<< polysilicon >>
rect 17 53 22 54
rect 17 50 18 53
rect 21 50 22 53
rect 17 49 22 50
rect 32 53 37 54
rect 32 50 33 53
rect 36 50 37 53
rect 32 49 37 50
rect 11 45 16 46
rect 11 42 12 45
rect 15 42 16 45
rect 11 41 16 42
rect 13 38 15 41
rect 20 38 22 49
rect 26 45 31 46
rect 26 42 27 45
rect 30 42 31 45
rect 26 41 31 42
rect 27 38 29 41
rect 34 38 36 49
rect 13 16 15 23
rect 20 16 22 23
rect 27 16 29 23
rect 34 16 36 23
rect 13 4 15 6
rect 20 4 22 6
rect 27 4 29 6
rect 34 4 36 6
<< pc >>
rect 18 50 21 53
rect 33 50 36 53
rect 12 42 15 45
rect 27 42 30 45
<< m1 >>
rect 3 13 6 58
rect 12 45 15 58
rect 18 53 21 58
rect 18 49 21 50
rect 12 41 15 42
rect 27 45 30 58
rect 33 53 36 58
rect 33 49 36 50
rect 27 41 30 42
rect 9 28 12 29
rect 36 28 39 29
rect 45 31 48 58
rect 9 24 12 25
rect 22 24 23 27
rect 26 24 27 27
rect 36 25 37 28
rect 40 25 41 28
rect 24 22 27 24
rect 15 16 18 17
rect 15 15 19 16
rect 15 12 16 15
rect 16 11 19 12
rect 9 10 12 11
rect 30 10 33 11
rect 22 7 23 10
rect 26 7 27 10
rect 9 5 12 7
rect 24 5 27 7
rect 30 6 33 7
rect 36 7 37 10
rect 40 7 41 10
rect 36 5 39 7
<< m2c >>
rect 9 29 12 32
rect 36 29 39 32
rect 45 28 48 31
rect 3 10 6 13
rect 15 17 18 20
rect 24 19 27 22
rect 30 11 33 14
rect 9 2 12 5
rect 24 2 27 5
rect 36 2 39 5
<< m2 >>
rect 8 32 13 33
rect 8 30 9 32
rect -8 29 9 30
rect 12 30 13 32
rect 35 32 40 33
rect 35 30 36 32
rect 12 29 36 30
rect 39 30 40 32
rect 44 31 49 32
rect 44 30 45 31
rect 39 29 45 30
rect -8 28 45 29
rect 48 30 49 31
rect 48 28 55 30
rect 44 27 49 28
rect 23 22 28 23
rect 14 20 19 21
rect 23 20 24 22
rect 14 17 15 20
rect 18 19 24 20
rect 27 19 28 22
rect 18 18 28 19
rect 18 17 19 18
rect 14 16 19 17
rect 29 14 34 15
rect 2 13 7 14
rect 2 12 3 13
rect -8 10 3 12
rect 6 12 7 13
rect 29 12 30 14
rect 6 11 30 12
rect 33 12 34 14
rect 33 11 55 12
rect 6 10 55 11
rect 2 9 7 10
rect 8 5 13 6
rect 8 2 9 5
rect 12 4 13 5
rect 23 5 28 6
rect 23 4 24 5
rect 12 2 24 4
rect 27 4 28 5
rect 35 5 40 6
rect 35 4 36 5
rect 27 2 36 4
rect 39 2 40 5
rect 8 1 13 2
rect 23 1 28 2
rect 35 1 40 2
<< labels >>
rlabel ndiffusion 37 7 37 7 3 #3
rlabel pdiffusion 37 24 37 24 3 Vdd
rlabel polysilicon 35 17 35 17 3 A
rlabel polysilicon 35 22 35 22 3 A
rlabel polysilicon 28 17 28 17 3 B
rlabel polysilicon 28 22 28 22 3 B
rlabel ndiffusion 23 7 23 7 3 #3
rlabel pdiffusion 23 24 23 24 3 Y
rlabel polysilicon 21 17 21 17 3 D
rlabel polysilicon 21 22 21 22 3 D
rlabel ndiffusion 16 7 16 7 3 Y
rlabel polysilicon 14 22 14 22 3 C
rlabel ndiffusion 9 7 9 7 3 #3
rlabel pdiffusion 9 24 9 24 3 Vdd
rlabel m2 30 2 33 4 1 #3
rlabel polysilicon 14 17 14 17 3 C
rlabel m2 22 18 24 20 1 Y
rlabel m1 12 56 15 58 4 C
rlabel m1 18 56 21 58 5 D
rlabel m1 27 56 30 58 5 B
rlabel m1 33 56 36 58 5 A
rlabel m2c 4 11 4 11 3 GND
rlabel m2 43 11 43 11 7 GND
rlabel m1 30 7 30 7 1 GND
rlabel m1 3 56 6 58 4 GND
rlabel m2 -2 28 -2 28 3 Vdd
rlabel m2 49 29 49 29 7 Vdd
rlabel m1 45 56 48 58 5 Vdd
<< end >>
