magic
tech sky130l
timestamp 1659179486
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 10 20 12
rect 15 7 16 10
rect 19 7 20 10
rect 15 6 20 7
rect 22 10 27 12
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
rect 29 10 34 12
rect 29 7 30 10
rect 33 7 34 10
rect 29 6 34 7
<< ndc >>
rect 9 7 12 10
rect 16 7 19 10
rect 23 7 26 10
rect 30 7 33 10
<< ntransistor >>
rect 13 6 15 12
rect 20 6 22 12
rect 27 6 29 12
<< pdiffusion >>
rect 8 36 13 37
rect 8 33 9 36
rect 12 33 13 36
rect 8 30 13 33
rect 8 27 9 30
rect 12 27 13 30
rect 8 24 13 27
rect 8 21 9 24
rect 12 21 13 24
rect 8 19 13 21
rect 15 19 20 37
rect 22 19 27 37
rect 29 36 34 37
rect 29 33 30 36
rect 33 33 34 36
rect 29 30 34 33
rect 29 27 30 30
rect 33 27 34 30
rect 29 24 34 27
rect 29 21 30 24
rect 33 21 34 24
rect 29 19 34 21
<< pdc >>
rect 9 33 12 36
rect 9 27 12 30
rect 9 21 12 24
rect 30 33 33 36
rect 30 27 33 30
rect 30 21 33 24
<< ptransistor >>
rect 13 19 15 37
rect 20 19 22 37
rect 27 19 29 37
<< polysilicon >>
rect 20 46 31 47
rect 20 43 21 46
rect 24 43 27 46
rect 30 43 31 46
rect 20 42 31 43
rect 13 37 15 39
rect 20 37 22 42
rect 27 37 29 39
rect 13 12 15 19
rect 20 12 22 19
rect 27 12 29 19
rect 13 1 15 6
rect 20 4 22 6
rect 27 1 29 6
rect 8 0 19 1
rect 8 -3 9 0
rect 12 -3 15 0
rect 18 -3 19 0
rect 8 -4 19 -3
rect 23 0 34 1
rect 23 -3 24 0
rect 27 -3 30 0
rect 33 -3 34 0
rect 23 -4 34 -3
<< pc >>
rect 21 43 24 46
rect 27 43 30 46
rect 9 -3 12 0
rect 15 -3 18 0
rect 24 -3 27 0
rect 30 -3 33 0
<< m1 >>
rect 20 43 21 46
rect 24 43 27 46
rect 30 43 31 46
rect 9 36 12 37
rect 9 30 12 33
rect 9 24 12 27
rect 9 20 12 21
rect 30 36 33 37
rect 30 30 33 33
rect 30 24 33 27
rect 30 18 33 21
rect 16 15 33 18
rect 9 10 12 11
rect 9 6 12 7
rect 16 10 19 15
rect 16 6 19 7
rect 23 10 26 11
rect 23 6 26 7
rect 30 10 33 15
rect 30 6 33 7
rect 8 -3 9 0
rect 12 -3 15 0
rect 18 -3 19 0
rect 23 -3 24 0
rect 27 -3 30 0
rect 33 -3 34 0
<< m2c >>
rect 9 33 12 36
rect 9 27 12 30
rect 9 7 12 10
rect 23 7 26 10
<< m2 >>
rect 8 36 13 37
rect 8 33 9 36
rect 12 33 13 36
rect 8 30 13 33
rect 8 27 9 30
rect 12 27 13 30
rect 8 26 13 27
rect 8 10 27 11
rect 8 7 9 10
rect 12 7 23 10
rect 26 7 27 10
rect 8 6 27 7
<< labels >>
rlabel ndiffusion 30 7 30 7 3 out
rlabel pdiffusion 30 20 30 20 3 out
rlabel polysilicon 28 13 28 13 3 in(2)
rlabel polysilicon 28 18 28 18 3 in(2)
rlabel ndiffusion 23 7 23 7 3 GND
rlabel polysilicon 21 13 21 13 3 in(1)
rlabel polysilicon 21 18 21 18 3 in(1)
rlabel ndiffusion 16 7 16 7 3 out
rlabel polysilicon 14 13 14 13 3 in(0)
rlabel polysilicon 14 18 14 18 3 in(0)
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 20 9 20 3 Vdd
flabel m2 8 26 13 37 0 FreeSans 11 0 0 0 Vdd
port 1 nsew
flabel m2 8 6 27 11 0 FreeSans 11 0 0 0 GND
flabel m1 8 -3 19 0 0 FreeSans 11 0 0 0 in(0)
port 3 nsew
flabel m1 20 43 31 46 0 FreeSans 11 0 0 0 in(1)
port 4 nsew
flabel m1 23 -3 34 0 0 FreeSans 11 0 0 0 in(2)
port 5 nsew
flabel m1 16 15 33 18 0 FreeSans 11 0 0 0 out
<< end >>
