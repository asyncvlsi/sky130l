magic
tech sky130l
timestamp 1636052260
<< ndiffusion >>
rect 6 15 11 16
rect 6 12 7 15
rect 10 12 11 15
rect 6 6 11 12
rect 13 6 18 16
rect 20 15 25 16
rect 20 12 21 15
rect 24 12 25 15
rect 20 10 25 12
rect 27 15 32 16
rect 27 12 28 15
rect 31 12 32 15
rect 27 10 32 12
rect 20 6 24 10
<< ndc >>
rect 7 12 10 15
rect 21 12 24 15
rect 28 12 31 15
<< ntransistor >>
rect 11 6 13 16
rect 18 6 20 16
rect 25 10 27 16
<< pdiffusion >>
rect 6 30 11 31
rect 6 27 7 30
rect 10 27 11 30
rect 6 23 11 27
rect 13 27 18 31
rect 13 24 14 27
rect 17 24 18 27
rect 13 23 18 24
rect 20 30 25 31
rect 20 27 21 30
rect 24 27 25 30
rect 20 23 25 27
rect 27 27 32 31
rect 27 24 28 27
rect 31 24 32 27
rect 27 23 32 24
<< pdc >>
rect 7 27 10 30
rect 14 24 17 27
rect 21 27 24 30
rect 28 24 31 27
<< ptransistor >>
rect 11 23 13 31
rect 18 23 20 31
rect 25 23 27 31
<< polysilicon >>
rect 8 38 13 39
rect 8 35 9 38
rect 12 35 13 38
rect 8 34 13 35
rect 17 38 22 39
rect 17 35 18 38
rect 21 35 22 38
rect 17 34 22 35
rect 11 31 13 34
rect 18 31 20 34
rect 25 31 27 33
rect 11 16 13 23
rect 18 16 20 23
rect 25 16 27 23
rect 11 4 13 6
rect 18 4 20 6
rect 25 5 27 10
rect 25 4 31 5
rect 25 3 27 4
rect 26 1 27 3
rect 30 1 31 4
rect 26 0 31 1
<< pc >>
rect 9 35 12 38
rect 18 35 21 38
rect 27 1 30 4
<< m1 >>
rect 9 38 12 42
rect 9 34 12 35
rect 18 38 21 42
rect 18 34 21 35
rect 6 30 11 31
rect 6 27 7 30
rect 10 27 11 30
rect 20 30 25 31
rect 6 26 11 27
rect 14 27 17 28
rect 20 27 21 30
rect 24 27 25 30
rect 20 26 25 27
rect 28 27 33 28
rect 14 23 17 24
rect 31 24 33 27
rect 28 23 33 24
rect 12 20 18 23
rect 12 16 15 20
rect 30 16 33 23
rect 6 15 15 16
rect 6 12 7 15
rect 10 12 15 15
rect 12 4 15 12
rect 20 15 25 16
rect 20 12 21 15
rect 24 12 25 15
rect 20 11 25 12
rect 28 15 33 16
rect 31 12 33 15
rect 28 11 33 12
rect 12 1 27 4
rect 30 1 31 4
rect 12 0 31 1
<< m2c >>
rect 7 27 10 30
rect 21 27 24 30
rect 21 12 24 15
<< m2 >>
rect 24 31 27 42
rect 6 30 11 31
rect 6 27 7 30
rect 10 28 11 30
rect 20 30 27 31
rect 20 28 21 30
rect 10 27 21 28
rect 24 28 27 30
rect 24 27 25 28
rect 6 26 25 27
rect 20 15 25 16
rect 20 12 21 15
rect 24 12 25 15
rect 20 10 25 12
rect 21 -2 24 10
<< labels >>
rlabel ndiffusion 28 11 28 11 3 Y
rlabel polysilicon 26 17 26 17 3 _Y
rlabel polysilicon 26 22 26 22 3 _Y
rlabel pdiffusion 28 24 28 24 3 Y
rlabel ndiffusion 21 7 21 7 3 GND
rlabel pdiffusion 21 24 21 24 3 Vdd
rlabel polysilicon 19 17 19 17 3 A
rlabel polysilicon 19 22 19 22 3 A
rlabel pdiffusion 14 24 14 24 3 _Y
rlabel polysilicon 12 17 12 17 3 B
rlabel polysilicon 12 22 12 22 3 B
rlabel ndiffusion 7 7 7 7 3 _Y
rlabel pdiffusion 7 24 7 24 3 Vdd
rlabel m1 31 19 31 19 3 Y
port 4 e
rlabel m1 10 40 10 40 3 B
port 3 e
rlabel m1 19 40 19 40 3 A
port 5 e
rlabel m2 25 41 25 41 3 Vdd
port 2 e
rlabel m2 22 -1 22 -1 3 GND
port 1 e
<< end >>
