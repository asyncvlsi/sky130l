magic
tech sky130l
timestamp 1636078168
<< ndiffusion >>
rect 8 15 13 16
rect 8 12 9 15
rect 12 12 13 15
rect 8 10 13 12
rect 41 10 44 16
rect 46 14 53 16
rect 46 11 48 14
rect 51 11 53 14
rect 46 10 53 11
rect 49 6 53 10
rect 55 6 58 16
rect 60 15 65 16
rect 60 12 61 15
rect 64 12 65 15
rect 60 10 65 12
rect 69 15 74 16
rect 69 12 70 15
rect 73 12 74 15
rect 69 10 74 12
rect 60 6 64 10
<< ndc >>
rect 9 12 12 15
rect 48 11 51 14
rect 61 12 64 15
rect 70 12 73 15
<< ntransistor >>
rect 13 10 41 16
rect 44 10 46 16
rect 53 6 55 16
rect 58 6 60 16
rect 65 10 69 16
<< pdiffusion >>
rect 49 29 53 35
rect 8 27 13 29
rect 8 24 9 27
rect 12 24 13 27
rect 8 23 13 24
rect 27 23 44 29
rect 46 28 53 29
rect 46 25 48 28
rect 51 25 53 28
rect 46 23 53 25
rect 55 23 58 35
rect 60 33 64 35
rect 60 27 65 33
rect 60 24 61 27
rect 64 24 65 27
rect 60 23 65 24
rect 69 27 74 33
rect 69 24 70 27
rect 73 24 74 27
rect 69 23 74 24
<< pdc >>
rect 9 24 12 27
rect 48 25 51 28
rect 61 24 64 27
rect 70 24 73 27
<< ptransistor >>
rect 13 23 27 29
rect 44 23 46 29
rect 53 23 55 35
rect 58 23 60 35
rect 65 23 69 33
<< polysilicon >>
rect 20 36 25 37
rect 20 33 21 36
rect 24 33 25 36
rect 20 31 25 33
rect 41 36 46 37
rect 41 33 42 36
rect 45 33 46 36
rect 53 35 55 37
rect 58 35 60 37
rect 41 32 46 33
rect 13 29 27 31
rect 44 29 46 32
rect 65 33 69 35
rect 13 21 27 23
rect 13 16 41 18
rect 44 16 46 23
rect 53 16 55 23
rect 58 16 60 23
rect 65 16 69 23
rect 13 8 41 10
rect 44 8 46 10
rect 35 7 40 8
rect 35 4 36 7
rect 39 4 40 7
rect 65 8 69 10
rect 66 7 71 8
rect 53 4 55 6
rect 35 3 40 4
rect 50 3 55 4
rect 50 0 51 3
rect 54 0 55 3
rect 50 -1 55 0
rect 58 4 60 6
rect 66 4 67 7
rect 70 4 71 7
rect 58 3 63 4
rect 66 3 71 4
rect 58 0 59 3
rect 62 0 63 3
rect 58 -1 63 0
<< pc >>
rect 21 33 24 36
rect 42 33 45 36
rect 36 4 39 7
rect 51 0 54 3
rect 67 4 70 7
rect 59 0 62 3
<< m1 >>
rect 21 36 24 37
rect 8 24 9 27
rect 12 24 13 27
rect 21 15 24 33
rect 42 36 45 37
rect 42 32 45 33
rect 48 28 51 29
rect 8 12 9 15
rect 12 12 13 15
rect 27 18 28 21
rect 27 7 30 18
rect 36 7 39 23
rect 72 27 75 33
rect 48 20 51 25
rect 60 24 61 27
rect 64 24 65 27
rect 69 24 70 27
rect 73 24 75 27
rect 48 14 51 17
rect 72 15 75 24
rect 60 12 61 15
rect 64 12 65 15
rect 69 12 70 15
rect 73 12 75 15
rect 72 11 75 12
rect 48 10 51 11
rect 66 4 67 7
rect 70 4 71 7
rect 36 3 39 4
rect 51 3 54 4
rect 51 -1 54 0
rect 59 3 62 4
rect 59 -1 62 0
rect 66 -1 69 4
<< m2c >>
rect 9 24 12 27
rect 42 33 45 36
rect 72 33 75 36
rect 36 23 39 26
rect 9 12 12 15
rect 21 12 24 15
rect 28 18 31 21
rect 27 4 30 7
rect 61 24 64 27
rect 48 17 51 20
rect 61 12 64 15
<< m2 >>
rect 41 36 46 37
rect 71 36 76 37
rect 41 33 42 36
rect 45 34 72 36
rect 45 33 46 34
rect 41 32 46 33
rect 71 33 72 34
rect 75 33 76 36
rect 71 32 76 33
rect 8 27 13 28
rect 60 27 65 28
rect 8 24 9 27
rect 12 26 13 27
rect 35 26 40 27
rect 60 26 61 27
rect 12 24 36 26
rect 8 23 13 24
rect 35 23 36 24
rect 39 24 61 26
rect 64 24 65 27
rect 39 23 40 24
rect 60 23 65 24
rect 35 22 40 23
rect 27 21 32 22
rect 27 18 28 21
rect 31 20 32 21
rect 47 20 52 21
rect 31 18 48 20
rect 27 17 32 18
rect 47 17 48 18
rect 51 17 52 20
rect 47 16 52 17
rect 8 15 13 16
rect 8 12 9 15
rect 12 14 13 15
rect 20 15 25 16
rect 20 14 21 15
rect 12 12 21 14
rect 24 14 25 15
rect 60 15 65 16
rect 60 14 61 15
rect 24 12 61 14
rect 64 12 65 15
rect 8 11 13 12
rect 20 11 25 12
rect 60 11 65 12
rect 26 7 31 8
rect 26 4 27 7
rect 30 6 31 7
rect 66 6 71 8
rect 30 4 71 6
rect 26 3 31 4
rect 66 3 71 4
<< labels >>
rlabel pdiffusion 70 24 70 24 3 #7
rlabel polysilicon 66 17 66 17 3 out
rlabel polysilicon 66 22 66 22 3 out
rlabel ndiffusion 70 11 70 11 3 #7
rlabel pdiffusion 61 24 61 24 3 Vdd
rlabel polysilicon 59 17 59 17 3 in(0)
rlabel polysilicon 59 22 59 22 3 in(0)
rlabel ndiffusion 61 7 61 7 3 GND
rlabel polysilicon 54 17 54 17 3 in(1)
rlabel polysilicon 54 22 54 22 3 in(1)
rlabel ndiffusion 47 11 47 11 3 out
rlabel pdiffusion 47 24 47 24 3 out
rlabel polysilicon 45 17 45 17 3 #7
rlabel polysilicon 45 22 45 22 3 #7
rlabel polysilicon 14 17 14 17 3 Vdd
rlabel polysilicon 14 22 14 22 3 GND
rlabel ndiffusion 9 11 9 11 3 GND
rlabel pdiffusion 9 24 9 24 3 Vdd
rlabel pc 53 1 53 1 3 in(1)
port 3 e
rlabel m2c 10 25 10 25 3 Vdd
port 2 e
rlabel pc 61 1 61 1 3 in(0)
port 5 e
rlabel m1 68 0 68 0 3 out
port 4 e
rlabel m1 9 13 9 13 3 GND
port 1 e
<< end >>
