magic
tech sky130l
timestamp 1639112566
<< ndiffusion >>
rect 8 10 13 16
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 15 20 16
rect 15 12 16 15
rect 19 12 20 15
rect 15 6 20 12
<< ndc >>
rect 9 7 12 10
rect 16 12 19 15
<< ntransistor >>
rect 13 6 15 16
<< pdiffusion >>
rect 8 27 13 38
rect 8 24 9 27
rect 12 24 13 27
rect 8 23 13 24
rect 15 27 20 38
rect 15 24 16 27
rect 19 24 20 27
rect 15 23 20 24
<< pdc >>
rect 9 24 12 27
rect 16 24 19 27
<< ptransistor >>
rect 13 23 15 38
<< polysilicon >>
rect 13 38 15 40
rect 13 16 15 23
rect 13 2 15 6
rect 11 1 16 2
rect 11 -2 12 1
rect 15 -2 16 1
rect 11 -3 16 -2
<< pc >>
rect 12 -2 15 1
<< m1 >>
rect 9 27 12 28
rect 9 23 12 24
rect 10 20 12 23
rect 15 27 21 28
rect 15 24 16 27
rect 19 24 21 27
rect 15 22 21 24
rect 15 16 18 22
rect 15 15 21 16
rect 15 12 16 15
rect 19 12 21 15
rect 9 10 12 12
rect 15 10 21 12
rect 6 9 9 10
rect 7 7 9 9
rect 7 6 12 7
rect 12 1 15 2
rect 12 -4 15 -2
<< m2c >>
rect 7 20 10 23
rect 4 6 7 9
<< m2 >>
rect 6 23 12 24
rect 6 22 7 23
rect 0 20 7 22
rect 10 20 12 23
rect 6 18 12 20
rect 3 9 9 10
rect 3 8 4 9
rect -3 6 4 8
rect 7 6 9 9
rect 3 4 9 6
<< labels >>
rlabel ndiffusion 16 7 16 7 3 out
rlabel pdiffusion 16 24 16 24 3 out
rlabel polysilicon 14 5 14 5 3 in(0)
rlabel ntransistor 14 7 14 7 3 in(0)
rlabel polysilicon 14 17 14 17 3 in(0)
rlabel polysilicon 14 22 14 22 3 in(0)
rlabel ptransistor 14 24 14 24 3 in(0)
rlabel polysilicon 14 39 14 39 3 in(0)
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 24 9 24 3 Vdd
rlabel m2 -3 6 0 8 2 GND
rlabel m2 0 20 3 22 3 Vdd
rlabel m1 12 -4 15 -3 1 in(0)
rlabel m1 15 18 18 20 7 out
<< end >>
