magic
tech sky130l
timestamp 1639255210
<< ndiffusion >>
rect 8 15 13 16
rect 8 12 9 15
rect 12 12 13 15
rect 8 10 13 12
rect 15 14 20 16
rect 15 11 16 14
rect 19 11 20 14
rect 15 10 20 11
rect 22 15 27 16
rect 22 12 23 15
rect 26 12 27 15
rect 22 10 27 12
rect 34 15 39 16
rect 34 12 35 15
rect 38 12 39 15
rect 34 6 39 12
rect 41 15 46 16
rect 41 12 42 15
rect 45 12 46 15
rect 41 6 46 12
rect 48 10 53 16
rect 48 7 49 10
rect 52 7 53 10
rect 48 6 53 7
rect 60 15 65 16
rect 60 12 61 15
rect 64 12 65 15
rect 60 6 65 12
rect 67 10 72 16
rect 67 7 68 10
rect 71 7 72 10
rect 67 6 72 7
rect 74 10 79 16
rect 74 7 75 10
rect 78 7 79 10
rect 74 6 79 7
<< ndc >>
rect 9 12 12 15
rect 16 11 19 14
rect 23 12 26 15
rect 35 12 38 15
rect 42 12 45 15
rect 49 7 52 10
rect 61 12 64 15
rect 68 7 71 10
rect 75 7 78 10
<< ntransistor >>
rect 13 10 15 16
rect 20 10 22 16
rect 39 6 41 16
rect 46 6 48 16
rect 65 6 67 16
rect 72 6 74 16
<< pdiffusion >>
rect 8 27 13 31
rect 8 24 9 27
rect 12 24 13 27
rect 8 23 13 24
rect 15 30 20 31
rect 15 27 16 30
rect 19 27 20 30
rect 15 23 20 27
rect 22 27 27 31
rect 22 24 23 27
rect 26 24 27 27
rect 22 23 27 24
rect 34 27 39 38
rect 34 24 35 27
rect 38 24 39 27
rect 34 23 39 24
rect 41 27 46 38
rect 41 24 42 27
rect 45 24 46 27
rect 41 23 46 24
rect 48 27 53 38
rect 48 24 49 27
rect 52 24 53 27
rect 48 23 53 24
rect 60 27 65 38
rect 60 24 61 27
rect 64 24 65 27
rect 60 23 65 24
rect 67 37 72 38
rect 67 34 68 37
rect 71 34 72 37
rect 67 23 72 34
rect 74 27 79 38
rect 74 24 75 27
rect 78 24 79 27
rect 74 23 79 24
<< pdc >>
rect 9 24 12 27
rect 16 27 19 30
rect 23 24 26 27
rect 35 24 38 27
rect 42 24 45 27
rect 49 24 52 27
rect 61 24 64 27
rect 68 34 71 37
rect 75 24 78 27
<< ptransistor >>
rect 13 23 15 31
rect 20 23 22 31
rect 39 23 41 38
rect 46 23 48 38
rect 65 23 67 38
rect 72 23 74 38
<< polysilicon >>
rect 8 45 15 46
rect 8 42 9 45
rect 12 42 15 45
rect 8 41 15 42
rect 36 45 41 46
rect 36 42 37 45
rect 40 42 41 45
rect 36 41 41 42
rect 13 31 15 41
rect 20 40 26 41
rect 20 37 22 40
rect 25 37 26 40
rect 39 38 41 41
rect 46 45 51 46
rect 46 42 47 45
rect 50 42 51 45
rect 46 41 51 42
rect 62 45 67 46
rect 62 42 63 45
rect 66 42 67 45
rect 74 45 79 46
rect 74 42 75 45
rect 78 42 79 45
rect 62 41 67 42
rect 46 38 48 41
rect 65 38 67 41
rect 72 41 79 42
rect 72 40 76 41
rect 72 38 74 40
rect 20 36 26 37
rect 20 31 22 36
rect 13 16 15 23
rect 20 16 22 23
rect 39 16 41 23
rect 46 16 48 23
rect 65 16 67 23
rect 72 16 74 23
rect 13 8 15 10
rect 20 8 22 10
rect 39 4 41 6
rect 46 4 48 6
rect 65 4 67 6
rect 72 4 74 6
<< pc >>
rect 9 42 12 45
rect 37 42 40 45
rect 22 37 25 40
rect 47 42 50 45
rect 63 42 66 45
rect 75 42 78 45
<< m1 >>
rect 8 45 12 46
rect 8 42 9 45
rect 8 41 12 42
rect 9 34 12 35
rect 9 27 12 31
rect 15 31 18 49
rect 36 45 42 46
rect 21 42 37 45
rect 40 42 42 45
rect 46 45 51 46
rect 46 42 47 45
rect 50 42 51 45
rect 21 40 25 42
rect 46 41 51 42
rect 63 45 66 46
rect 63 41 66 42
rect 21 37 22 40
rect 21 36 25 37
rect 48 35 51 41
rect 69 38 72 49
rect 35 34 51 35
rect 29 33 51 34
rect 68 37 72 38
rect 71 34 72 37
rect 68 33 72 34
rect 75 45 78 46
rect 75 34 78 42
rect 23 32 51 33
rect 23 31 38 32
rect 15 30 19 31
rect 15 27 16 30
rect 15 26 19 27
rect 23 30 32 31
rect 23 27 26 30
rect 9 15 12 24
rect 23 15 26 24
rect 35 27 39 28
rect 38 24 39 27
rect 35 23 39 24
rect 42 27 45 28
rect 75 27 78 28
rect 48 24 49 27
rect 52 24 61 27
rect 64 24 65 27
rect 78 24 79 27
rect 9 11 12 12
rect 15 14 19 15
rect 15 11 16 14
rect 23 11 26 12
rect 35 15 39 16
rect 38 12 39 15
rect 35 11 39 12
rect 42 15 45 24
rect 75 23 78 24
rect 15 10 19 11
rect 15 2 18 10
rect 42 4 45 12
rect 60 15 64 16
rect 60 12 61 15
rect 60 11 64 12
rect 48 10 52 11
rect 48 7 49 10
rect 48 6 52 7
rect 68 10 72 11
rect 71 7 72 10
rect 68 6 72 7
rect 75 10 78 11
rect 75 6 78 7
rect 69 2 72 6
rect 15 -2 18 -1
<< m2c >>
rect 15 49 18 52
rect 9 42 12 45
rect 9 31 12 34
rect 69 49 72 52
rect 63 42 66 45
rect 75 31 78 34
rect 35 24 38 27
rect 79 24 82 27
rect 35 12 38 15
rect 61 12 64 15
rect 49 7 52 10
rect 75 7 78 10
rect 15 -1 18 2
rect 69 -1 72 2
<< m2 >>
rect 14 52 73 53
rect 14 49 15 52
rect 18 49 69 52
rect 72 49 73 52
rect 14 48 73 49
rect 8 45 67 46
rect 8 42 9 45
rect 12 44 63 45
rect 12 42 13 44
rect 8 41 13 42
rect 62 42 63 44
rect 66 42 67 45
rect 62 41 67 42
rect 8 34 13 35
rect 8 31 9 34
rect 12 32 13 34
rect 74 34 79 35
rect 74 32 75 34
rect 12 31 75 32
rect 78 31 79 34
rect 8 30 79 31
rect 34 27 39 28
rect 34 24 35 27
rect 38 26 39 27
rect 78 27 83 28
rect 78 26 79 27
rect 38 24 79 26
rect 82 24 83 27
rect 34 23 39 24
rect 78 23 83 24
rect 34 15 65 16
rect 34 12 35 15
rect 38 14 61 15
rect 38 12 39 14
rect 34 11 39 12
rect 60 12 61 14
rect 64 12 65 15
rect 60 11 65 12
rect 48 10 53 11
rect 48 7 49 10
rect 52 8 53 10
rect 74 10 79 11
rect 74 8 75 10
rect 52 7 75 8
rect 78 7 79 10
rect 48 6 79 7
rect 14 2 73 3
rect 14 -1 15 2
rect 18 -1 69 2
rect 72 -1 73 2
rect 14 -2 73 -1
<< labels >>
rlabel ndiffusion 61 7 61 7 3 #10
rlabel pdiffusion 68 24 68 24 3 Vdd
rlabel pdiffusion 42 24 42 24 3 Y
rlabel ndiffusion 42 7 42 7 3 Y
rlabel pdiffusion 49 24 49 24 3 #7
rlabel pdiffusion 9 24 9 24 3 _B
rlabel ndiffusion 9 11 9 11 3 _B
rlabel polysilicon 14 17 14 17 3 B
rlabel pdiffusion 16 24 16 24 3 Vdd
rlabel ndiffusion 16 11 16 11 3 GND
rlabel polysilicon 21 17 21 17 3 A
rlabel pdiffusion 23 24 23 24 3 _A
rlabel ndiffusion 23 11 23 11 3 _A
rlabel ndiffusion 35 7 35 7 1 #10
rlabel pdiffusion 62 30 62 30 1 #7
rlabel pdiffusion 75 30 75 30 1 #8
rlabel polysilicon 66 22 66 22 1 B
rlabel polysilicon 66 17 66 17 1 B
rlabel polysilicon 73 22 73 22 1 _B
rlabel polysilicon 73 17 73 17 1 _B
rlabel polysilicon 40 22 40 22 1 A
rlabel polysilicon 40 17 40 17 1 A
rlabel polysilicon 47 22 47 22 1 _A
rlabel polysilicon 47 17 47 17 1 _A
rlabel m1 37 43 37 43 3 A
port 5 e
rlabel ndiffusion 76 7 76 7 3 #9
rlabel ndiffusion 50 7 50 7 1 #9
rlabel m1 70 10 70 10 1 GND
rlabel m1 43 5 43 5 3 Y
port 4 e
rlabel m2c 71 0 71 0 1 GND
rlabel m1 16 -1 16 -1 3 GND
port 1 e
rlabel m2c 62 14 62 14 1 #10
rlabel m2c 16 50 16 50 3 Vdd
port 2 e
rlabel m2c 71 50 71 50 5 Vdd
rlabel polysilicon 21 22 21 22 3 A
rlabel polysilicon 14 22 14 22 3 B
<< end >>
