magic
tech sky130l
timestamp 1636602381
<< ndiffusion >>
rect 6 12 11 16
rect 6 9 7 12
rect 10 9 11 12
rect 6 6 11 9
rect 13 6 18 16
rect 20 15 25 16
rect 20 12 21 15
rect 24 12 25 15
rect 20 10 25 12
rect 27 14 32 16
rect 27 11 28 14
rect 31 11 32 14
rect 27 10 32 11
rect 20 6 24 10
<< ndc >>
rect 7 9 10 12
rect 21 12 24 15
rect 28 11 31 14
<< ntransistor >>
rect 11 6 13 16
rect 18 6 20 16
rect 25 10 27 16
<< pdiffusion >>
rect 6 35 11 38
rect 6 32 7 35
rect 10 32 11 35
rect 6 23 11 32
rect 13 27 18 38
rect 13 24 14 27
rect 17 24 18 27
rect 13 23 18 24
rect 20 35 25 38
rect 20 32 21 35
rect 24 32 25 35
rect 20 23 25 32
rect 27 27 32 38
rect 27 24 28 27
rect 31 24 32 27
rect 27 23 32 24
<< pdc >>
rect 7 32 10 35
rect 14 24 17 27
rect 21 32 24 35
rect 28 24 31 27
<< ptransistor >>
rect 11 23 13 38
rect 18 23 20 38
rect 25 23 27 38
<< polysilicon >>
rect 8 45 13 46
rect 8 42 9 45
rect 12 42 13 45
rect 8 41 13 42
rect 17 45 22 46
rect 17 42 18 45
rect 21 42 22 45
rect 26 45 31 46
rect 26 43 27 45
rect 17 41 22 42
rect 25 42 27 43
rect 30 42 31 45
rect 25 41 31 42
rect 11 38 13 41
rect 18 38 20 41
rect 25 38 27 41
rect 11 16 13 23
rect 18 16 20 23
rect 25 16 27 23
rect 25 8 27 10
rect 11 4 13 6
rect 18 4 20 6
<< pc >>
rect 9 42 12 45
rect 18 42 21 45
rect 27 42 30 45
<< m1 >>
rect 9 45 12 49
rect 9 41 12 42
rect 18 45 21 49
rect 18 41 21 42
rect 27 45 30 49
rect 27 41 30 42
rect 6 35 25 36
rect 6 32 7 35
rect 10 32 21 35
rect 24 32 25 35
rect 13 27 18 28
rect 13 24 14 27
rect 17 24 18 27
rect 13 23 18 24
rect 27 24 28 27
rect 31 24 32 27
rect 27 22 30 24
rect 21 18 30 22
rect 21 15 24 18
rect 6 12 11 13
rect 6 9 7 12
rect 10 9 11 12
rect 6 8 11 9
rect 21 2 24 12
rect 27 14 32 15
rect 27 11 28 14
rect 31 11 32 14
rect 27 10 32 11
<< m2c >>
rect 14 24 17 27
rect 7 9 10 12
rect 28 11 31 14
<< m2 >>
rect 13 27 18 28
rect 13 26 14 27
rect -9 24 14 26
rect 17 24 18 27
rect 13 23 18 24
rect 27 14 32 15
rect 6 12 11 13
rect 27 12 28 14
rect 3 10 7 12
rect 6 9 7 10
rect 10 11 28 12
rect 31 11 32 14
rect 10 10 32 11
rect 10 9 11 10
rect 6 8 11 9
<< labels >>
rlabel ndiffusion 28 11 28 11 3 GND
rlabel polysilicon 26 17 26 17 3 C
rlabel polysilicon 26 22 26 22 3 C
rlabel pdiffusion 28 24 28 24 3 Y
rlabel ndiffusion 21 7 21 7 3 Y
rlabel pdiffusion 21 24 21 24 3 #7
rlabel polysilicon 19 17 19 17 3 B
rlabel polysilicon 19 22 19 22 3 B
rlabel pdiffusion 14 24 14 24 3 Vdd
rlabel polysilicon 12 17 12 17 3 A
rlabel polysilicon 12 22 12 22 3 A
rlabel pdiffusion 7 24 7 24 3 #7
rlabel ndiffusion 7 7 7 7 3 GND
rlabel m1 10 47 10 47 3 A
port 6 e
rlabel m1 19 47 19 47 3 B
port 4 e
rlabel m1 28 47 28 47 3 C
port 3 e
rlabel m2 4 25 4 25 3 Vdd
port 2 e
rlabel m2 4 11 4 11 3 GND
port 1 e
rlabel m1 22 3 22 3 3 Y
port 5 e
<< end >>
