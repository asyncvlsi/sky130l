magic
tech sky130l
timestamp 1659174961
<< ndiffusion >>
rect 8 12 13 16
rect 8 9 9 12
rect 12 9 13 12
rect 8 6 13 9
rect 15 12 20 16
rect 15 9 16 12
rect 19 9 20 12
rect 15 6 20 9
rect 22 6 27 16
rect 29 12 34 16
rect 29 9 30 12
rect 33 9 34 12
rect 29 6 34 9
rect 36 12 41 16
rect 36 9 37 12
rect 40 9 41 12
rect 36 6 41 9
rect 47 12 52 14
rect 47 9 48 12
rect 51 9 52 12
rect 47 8 52 9
rect 54 8 59 14
rect 87 12 92 14
rect 87 9 88 12
rect 91 9 92 12
rect 87 8 92 9
rect 96 12 102 14
rect 96 9 98 12
rect 101 9 102 12
rect 96 8 102 9
<< ndc >>
rect 9 9 12 12
rect 16 9 19 12
rect 30 9 33 12
rect 37 9 40 12
rect 48 9 51 12
rect 88 9 91 12
rect 98 9 101 12
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
rect 27 6 29 16
rect 34 6 36 16
rect 52 8 54 14
rect 59 8 87 14
rect 92 8 96 14
<< pdiffusion >>
rect 8 34 13 35
rect 8 31 9 34
rect 12 31 13 34
rect 8 28 13 31
rect 8 25 9 28
rect 12 25 13 28
rect 8 23 13 25
rect 15 23 20 35
rect 22 34 27 35
rect 22 31 23 34
rect 26 31 27 34
rect 87 31 92 35
rect 22 28 27 31
rect 47 30 52 31
rect 22 25 23 28
rect 26 25 27 28
rect 22 23 27 25
rect 47 27 48 30
rect 51 27 52 30
rect 47 25 52 27
rect 54 25 66 31
rect 80 30 92 31
rect 80 27 82 30
rect 85 27 88 30
rect 91 27 92 30
rect 80 25 92 27
rect 96 30 102 35
rect 96 27 98 30
rect 101 27 102 30
rect 96 25 102 27
<< pdc >>
rect 9 31 12 34
rect 9 25 12 28
rect 23 31 26 34
rect 23 25 26 28
rect 48 27 51 30
rect 82 27 85 30
rect 88 27 91 30
rect 98 27 101 30
<< ptransistor >>
rect 13 23 15 35
rect 20 23 22 35
rect 52 25 54 31
rect 66 25 80 31
rect 92 25 96 35
<< polysilicon >>
rect 20 42 31 43
rect 20 39 21 42
rect 24 39 27 42
rect 30 39 31 42
rect 20 38 31 39
rect 66 38 80 39
rect 13 35 15 37
rect 20 35 22 38
rect 66 35 67 38
rect 70 35 73 38
rect 76 35 80 38
rect 92 35 96 37
rect 52 31 54 33
rect 66 31 80 35
rect 32 27 43 28
rect 32 24 33 27
rect 36 24 39 27
rect 42 24 43 27
rect 32 23 43 24
rect 13 16 15 23
rect 20 16 22 23
rect 27 16 29 18
rect 34 16 36 23
rect 52 14 54 25
rect 66 23 80 25
rect 92 22 96 25
rect 90 21 96 22
rect 90 18 91 21
rect 94 18 96 21
rect 90 17 96 18
rect 59 14 87 16
rect 92 14 96 17
rect 13 0 15 6
rect 20 4 22 6
rect 27 0 29 6
rect 34 4 36 6
rect 52 0 54 8
rect 59 5 87 8
rect 92 6 96 8
rect 59 2 60 5
rect 63 2 66 5
rect 69 2 72 5
rect 75 2 78 5
rect 81 2 87 5
rect 59 1 87 2
rect 8 -1 19 0
rect 8 -4 9 -1
rect 12 -4 15 -1
rect 18 -4 19 -1
rect 8 -5 19 -4
rect 27 -1 38 0
rect 27 -4 28 -1
rect 31 -4 34 -1
rect 37 -4 38 -1
rect 27 -5 38 -4
rect 43 -1 54 0
rect 43 -4 44 -1
rect 47 -4 50 -1
rect 53 -4 54 -1
rect 43 -5 54 -4
<< pc >>
rect 21 39 24 42
rect 27 39 30 42
rect 67 35 70 38
rect 73 35 76 38
rect 33 24 36 27
rect 39 24 42 27
rect 91 18 94 21
rect 60 2 63 5
rect 66 2 69 5
rect 72 2 75 5
rect 78 2 81 5
rect 9 -4 12 -1
rect 15 -4 18 -1
rect 28 -4 31 -1
rect 34 -4 37 -1
rect 44 -4 47 -1
rect 50 -4 53 -1
<< m1 >>
rect 20 39 21 42
rect 24 39 27 42
rect 30 39 31 42
rect 57 35 67 38
rect 70 35 73 38
rect 76 35 77 38
rect 9 34 12 35
rect 9 28 12 31
rect 9 24 12 25
rect 23 34 26 35
rect 23 28 26 31
rect 48 30 51 31
rect 23 21 26 25
rect 32 24 33 27
rect 36 24 39 27
rect 42 24 43 27
rect 48 21 51 27
rect 57 27 62 35
rect 98 30 101 31
rect 81 27 82 30
rect 85 27 88 30
rect 91 27 92 30
rect 57 24 58 27
rect 61 24 62 27
rect 23 18 91 21
rect 94 18 95 21
rect 9 12 12 13
rect 9 5 12 9
rect 16 12 19 13
rect 16 8 19 9
rect 30 12 33 18
rect 30 8 33 9
rect 37 12 40 13
rect 37 5 40 9
rect 48 12 51 18
rect 48 8 51 9
rect 74 12 75 15
rect 78 12 81 15
rect 84 12 85 15
rect 88 12 91 13
rect 74 5 82 12
rect 88 8 91 9
rect 98 12 101 27
rect 9 2 40 5
rect 59 2 60 5
rect 63 2 66 5
rect 69 2 72 5
rect 75 2 78 5
rect 81 2 82 5
rect 98 -1 101 9
rect 8 -4 9 -1
rect 12 -4 15 -1
rect 18 -4 19 -1
rect 27 -4 28 -1
rect 31 -4 34 -1
rect 37 -4 38 -1
rect 43 -4 44 -1
rect 47 -4 50 -1
rect 53 -4 101 -1
<< m2c >>
rect 58 24 61 27
rect 75 12 78 15
rect 81 12 84 15
<< m2 >>
rect 8 33 13 35
rect 8 30 92 33
rect 8 24 13 30
rect 57 27 62 28
rect 57 24 58 27
rect 61 24 62 27
rect 15 9 20 13
rect 57 9 62 24
rect 74 26 92 30
rect 74 15 85 26
rect 74 12 75 15
rect 78 12 81 15
rect 84 12 85 15
rect 74 11 85 12
rect 87 9 92 13
rect 15 6 92 9
<< labels >>
rlabel ndiffusion 12 7 12 7 7 #3
rlabel pdiffusion 12 24 12 24 7 Vdd
rlabel polysilicon 14 17 14 17 7 in(0)
rlabel polysilicon 14 22 14 22 7 in(0)
rlabel ndiffusion 19 7 19 7 7 GND
rlabel polysilicon 21 17 21 17 7 in(2)
rlabel polysilicon 21 22 21 22 7 in(2)
rlabel pdiffusion 26 24 26 24 7 out
rlabel polysilicon 28 17 28 17 7 in(3)
rlabel ndiffusion 33 7 33 7 7 out
rlabel polysilicon 35 17 35 17 7 in(1)
rlabel ndiffusion 40 7 40 7 7 #3
rlabel pdiffusion 91 26 91 26 7 Vdd
rlabel polysilicon 95 24 95 24 7 out
rlabel pdiffusion 51 26 51 26 7 #11
rlabel polysilicon 53 24 53 24 7 #10
rlabel pdiffusion 58 26 58 26 7 out
rlabel pdiffusion 65 26 65 26 7 #11
rlabel polysilicon 79 24 79 24 7 GND
rlabel ndiffusion 48 9 48 9 3 out
rlabel polysilicon 53 15 53 15 3 #10
rlabel ndiffusion 55 9 55 9 3 #12
rlabel polysilicon 60 15 60 15 3 Vdd
rlabel ndiffusion 88 9 88 9 3 GND
rlabel polysilicon 93 15 93 15 3 out
rlabel pdiffusion 101 26 101 26 7 #10
rlabel ndiffusion 98 9 98 9 3 #10
flabel m2 8 30 92 33 0 FreeSans 11 0 0 0 Vdd
port 1 nsew
flabel m2 15 6 92 9 0 FreeSans 11 0 0 0 GND
flabel m1 8 -4 19 -1 0 FreeSans 11 0 0 0 in(0)
port 3 nsew
flabel m1 32 24 43 27 0 FreeSans 11 0 0 0 in(1)
port 4 nsew
flabel m1 20 39 31 42 0 FreeSans 11 0 0 0 in(2)
port 5 nsew
flabel m1 27 -4 38 -1 0 FreeSans 11 0 0 0 in(3)
port 6 nsew
flabel m1 23 18 95 21 0 FreeSans 11 0 0 0 out
port 7 nsew
<< end >>
