magic
tech sky130l
timestamp 1636155774
<< ndiffusion >>
rect 6 10 11 12
rect 6 7 7 10
rect 10 7 11 10
rect 6 6 11 7
rect 39 10 44 12
rect 39 7 40 10
rect 43 7 44 10
rect 39 6 44 7
rect 46 10 51 12
rect 46 7 47 10
rect 50 7 51 10
rect 46 6 51 7
rect 53 10 58 12
rect 53 7 54 10
rect 57 7 58 10
rect 53 6 58 7
rect 62 10 67 12
rect 62 7 63 10
rect 66 7 67 10
rect 62 6 67 7
rect 73 11 78 12
rect 73 8 74 11
rect 77 8 78 11
rect 73 6 78 8
rect 80 10 85 12
rect 80 7 81 10
rect 84 7 85 10
rect 80 6 85 7
<< ndc >>
rect 7 7 10 10
rect 40 7 43 10
rect 47 7 50 10
rect 54 7 57 10
rect 63 7 66 10
rect 74 8 77 11
rect 81 7 84 10
<< ntransistor >>
rect 11 6 39 12
rect 44 6 46 12
rect 51 6 53 12
rect 58 6 62 12
rect 78 6 80 12
<< pdiffusion >>
rect 6 23 11 37
rect 6 20 7 23
rect 10 20 11 23
rect 6 19 11 20
rect 13 19 44 37
rect 46 19 51 37
rect 53 29 57 37
rect 53 23 58 29
rect 53 20 54 23
rect 57 20 58 23
rect 53 19 58 20
rect 62 23 67 29
rect 62 20 63 23
rect 66 20 67 23
rect 62 19 67 20
rect 73 23 78 25
rect 73 20 74 23
rect 77 20 78 23
rect 73 19 78 20
rect 80 19 83 25
rect 94 23 99 25
rect 94 20 95 23
rect 98 20 99 23
rect 94 19 99 20
<< pdc >>
rect 7 20 10 23
rect 54 20 57 23
rect 63 20 66 23
rect 74 20 77 23
rect 95 20 98 23
<< ptransistor >>
rect 11 19 13 37
rect 44 19 46 37
rect 51 19 53 37
rect 58 19 62 29
rect 78 19 80 25
rect 83 19 94 25
<< polysilicon >>
rect 11 44 16 45
rect 11 41 12 44
rect 15 41 16 44
rect 11 40 16 41
rect 41 44 46 45
rect 41 41 42 44
rect 45 41 46 44
rect 41 40 46 41
rect 11 37 13 40
rect 44 37 46 40
rect 51 44 56 45
rect 51 41 52 44
rect 55 41 56 44
rect 51 40 56 41
rect 51 37 53 40
rect 75 32 80 33
rect 58 29 62 31
rect 75 29 76 32
rect 79 29 80 32
rect 75 28 80 29
rect 78 25 80 28
rect 83 25 94 27
rect 11 17 13 19
rect 11 12 39 14
rect 44 12 46 19
rect 51 12 53 19
rect 58 12 62 19
rect 78 12 80 19
rect 83 17 94 19
rect 89 15 94 17
rect 89 12 90 15
rect 93 12 94 15
rect 89 11 94 12
rect 11 4 39 6
rect 44 4 46 6
rect 51 4 53 6
rect 58 4 62 6
rect 78 4 80 6
rect 34 3 39 4
rect 34 0 35 3
rect 38 0 39 3
rect 34 -1 39 0
rect 57 3 62 4
rect 57 0 58 3
rect 61 0 62 3
rect 57 -1 62 0
<< pc >>
rect 12 41 15 44
rect 42 41 45 44
rect 52 41 55 44
rect 76 29 79 32
rect 90 12 93 15
rect 35 0 38 3
rect 58 0 61 3
<< m1 >>
rect 11 44 16 45
rect 41 44 46 45
rect 11 41 12 44
rect 15 41 16 44
rect 11 40 16 41
rect 9 24 12 25
rect 7 23 12 24
rect 10 20 12 23
rect 7 19 12 20
rect 9 17 12 19
rect 15 10 18 34
rect 6 7 7 10
rect 10 7 11 10
rect 33 23 36 41
rect 41 41 42 44
rect 45 41 46 44
rect 41 40 46 41
rect 51 44 56 45
rect 51 41 52 44
rect 55 41 56 44
rect 51 40 56 41
rect 63 32 66 33
rect 33 4 36 20
rect 47 10 50 25
rect 63 23 66 29
rect 76 32 79 33
rect 76 28 79 29
rect 74 23 77 24
rect 53 20 54 23
rect 57 20 58 23
rect 63 10 66 20
rect 39 7 40 10
rect 43 7 44 10
rect 53 7 54 10
rect 57 7 58 10
rect 33 3 39 4
rect 33 0 35 3
rect 38 0 39 3
rect 47 3 50 7
rect 63 6 66 7
rect 72 20 74 23
rect 72 19 77 20
rect 72 17 75 19
rect 72 12 75 14
rect 72 11 77 12
rect 72 8 74 11
rect 72 7 77 8
rect 80 7 81 10
rect 84 7 87 34
rect 96 23 99 41
rect 94 20 95 23
rect 98 20 99 23
rect 90 15 93 16
rect 90 10 93 12
rect 57 0 58 3
rect 61 0 62 3
rect 33 -1 39 0
rect 72 -1 75 7
rect 90 -1 93 7
<< m2c >>
rect 33 41 36 44
rect 15 34 18 37
rect 9 25 12 28
rect 9 14 12 17
rect 7 7 10 10
rect 15 7 18 10
rect 96 41 99 44
rect 84 34 87 37
rect 63 29 66 32
rect 33 20 36 23
rect 47 25 50 28
rect 76 29 79 32
rect 54 20 57 23
rect 40 7 43 10
rect 54 7 57 10
rect 72 14 75 17
rect 90 7 93 10
rect 47 0 50 3
rect 58 0 61 3
<< m2 >>
rect 32 44 37 45
rect 32 41 33 44
rect 36 42 37 44
rect 95 44 100 45
rect 95 42 96 44
rect 36 41 96 42
rect 99 41 100 44
rect 32 40 100 41
rect 14 37 88 38
rect 14 34 15 37
rect 18 36 84 37
rect 18 34 19 36
rect 14 33 19 34
rect 83 34 84 36
rect 87 34 88 37
rect 83 33 88 34
rect 62 32 67 33
rect 75 32 80 33
rect 62 29 63 32
rect 66 30 76 32
rect 66 29 67 30
rect 8 28 13 29
rect 46 28 51 29
rect 62 28 67 29
rect 75 29 76 30
rect 79 29 80 32
rect 75 28 80 29
rect 8 25 9 28
rect 12 26 47 28
rect 12 25 13 26
rect 8 24 13 25
rect 46 25 47 26
rect 50 25 51 28
rect 46 24 51 25
rect 32 23 37 24
rect 32 20 33 23
rect 36 22 37 23
rect 53 23 58 24
rect 53 22 54 23
rect 36 20 54 22
rect 57 20 58 23
rect 32 19 37 20
rect 53 19 58 20
rect 8 17 13 18
rect 8 14 9 17
rect 12 16 13 17
rect 71 17 76 18
rect 71 16 72 17
rect 12 14 72 16
rect 75 14 76 17
rect 8 13 13 14
rect 71 13 76 14
rect 6 10 11 11
rect 14 10 19 11
rect 6 7 7 10
rect 10 8 15 10
rect 10 7 11 8
rect 6 6 11 7
rect 14 7 15 8
rect 18 7 19 10
rect 14 6 19 7
rect 39 10 44 11
rect 39 7 40 10
rect 43 8 44 10
rect 53 10 58 11
rect 53 8 54 10
rect 43 7 54 8
rect 57 8 58 10
rect 89 10 94 11
rect 89 8 90 10
rect 57 7 90 8
rect 93 7 94 10
rect 39 6 94 7
rect 46 3 51 4
rect 46 0 47 3
rect 50 2 51 3
rect 57 3 62 4
rect 57 2 58 3
rect 50 0 58 2
rect 61 0 62 3
rect 46 -1 51 0
rect 57 -1 62 0
<< labels >>
rlabel pdiffusion 63 20 63 20 3 #8
rlabel ndiffusion 63 7 63 7 3 #8
rlabel polysilicon 59 13 59 13 3 out
rlabel polysilicon 59 18 59 18 3 out
rlabel ndiffusion 54 7 54 7 3 GND
rlabel pdiffusion 54 20 54 20 3 Vdd
rlabel polysilicon 52 13 52 13 3 in(0)
rlabel polysilicon 52 18 52 18 3 in(0)
rlabel ndiffusion 47 7 47 7 3 out
rlabel polysilicon 45 13 45 13 3 in(1)
rlabel polysilicon 45 18 45 18 3 in(1)
rlabel ndiffusion 40 7 40 7 3 GND
rlabel polysilicon 12 13 12 13 3 Vdd
rlabel polysilicon 12 18 12 18 3 in(2)
rlabel ndiffusion 7 7 7 7 3 #10
rlabel pdiffusion 7 20 7 20 3 out
rlabel pdiffusion 95 20 95 20 3 Vdd
rlabel polysilicon 84 18 84 18 3 GND
rlabel ndiffusion 81 7 81 7 3 #10
rlabel polysilicon 79 13 79 13 3 #8
rlabel polysilicon 79 18 79 18 3 #8
rlabel ndiffusion 74 7 74 7 3 out
rlabel pdiffusion 74 20 74 20 3 out
rlabel m1 74 1 74 1 3 out
port 5 e
rlabel pc 13 42 13 42 3 in(2)
port 3 e
rlabel m2c 35 42 35 42 3 Vdd
port 2 e
rlabel m1 92 1 92 1 3 GND
port 1 e
rlabel pc 44 44 44 44 3 in(1)
port 4 e
rlabel m1 55 44 55 44 3 in(0)
port 6 e
<< end >>
