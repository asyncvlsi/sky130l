magic
tech sky130l
timestamp 1659178732
<< ndiffusion >>
rect 8 12 13 16
rect 8 9 9 12
rect 12 9 13 12
rect 8 6 13 9
rect 15 6 20 16
rect 22 12 27 16
rect 22 9 23 12
rect 26 9 27 12
rect 22 6 27 9
<< ndc >>
rect 9 9 12 12
rect 23 9 26 12
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
<< pdiffusion >>
rect 8 28 13 29
rect 8 25 9 28
rect 12 25 13 28
rect 8 23 13 25
rect 15 28 20 29
rect 15 25 16 28
rect 19 25 20 28
rect 15 23 20 25
rect 22 28 27 29
rect 22 25 23 28
rect 26 25 27 28
rect 22 23 27 25
<< pdc >>
rect 9 25 12 28
rect 16 25 19 28
rect 23 25 26 28
<< ptransistor >>
rect 13 23 15 29
rect 20 23 22 29
<< polysilicon >>
rect 6 36 17 37
rect 6 33 7 36
rect 10 33 13 36
rect 16 33 17 36
rect 6 32 17 33
rect 13 29 15 32
rect 20 29 22 31
rect 13 16 15 23
rect 20 16 22 23
rect 13 4 15 6
rect 20 3 22 6
rect 18 2 29 3
rect 18 -1 19 2
rect 22 -1 25 2
rect 28 -1 29 2
rect 18 -2 29 -1
<< pc >>
rect 7 33 10 36
rect 13 33 16 36
rect 19 -1 22 2
rect 25 -1 28 2
<< m1 >>
rect 6 33 7 36
rect 10 33 13 36
rect 16 33 17 36
rect 9 28 12 29
rect 9 24 12 25
rect 16 28 19 29
rect 16 20 19 25
rect 23 28 26 29
rect 23 24 26 25
rect 16 17 26 20
rect 9 12 12 13
rect 9 8 12 9
rect 23 12 26 17
rect 23 8 26 9
rect 18 -1 19 2
rect 22 -1 25 2
rect 28 -1 29 2
<< m2c >>
rect 9 25 12 28
rect 23 25 26 28
rect 9 9 12 12
<< m2 >>
rect 8 28 27 29
rect 8 25 9 28
rect 12 25 23 28
rect 26 25 27 28
rect 8 24 27 25
rect 8 12 20 13
rect 8 9 9 12
rect 12 9 20 12
rect 8 8 20 9
<< labels >>
rlabel ndiffusion 23 7 23 7 3 out
rlabel pdiffusion 23 24 23 24 3 Vdd
rlabel polysilicon 21 17 21 17 3 in(1)
rlabel polysilicon 21 22 21 22 3 in(1)
rlabel pdiffusion 16 24 16 24 3 out
rlabel polysilicon 14 17 14 17 3 in(0)
rlabel polysilicon 14 22 14 22 3 in(0)
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 24 9 24 3 Vdd
flabel m2 8 24 27 29 0 FreeSans 11 0 0 0 Vdd
flabel m2 8 8 20 13 0 FreeSans 11 0 0 0 GND
port 2 nsew
flabel m1 6 33 17 36 0 FreeSans 11 0 0 0 in(0)
port 3 nsew
flabel m1 18 -1 29 2 0 FreeSans 11 0 0 0 in(1)
port 4 nsew
flabel m1 16 17 26 20 0 FreeSans 11 0 0 0 out
<< end >>
