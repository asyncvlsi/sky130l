magic
tech sky130l
timestamp 1659185046
<< ndiffusion >>
rect 8 9 13 12
rect 8 6 9 9
rect 12 6 13 9
rect 8 4 13 6
rect 15 9 20 12
rect 15 6 16 9
rect 19 6 20 9
rect 15 4 20 6
rect 22 9 27 12
rect 22 6 23 9
rect 26 6 27 9
rect 22 4 27 6
rect 29 9 34 12
rect 29 6 30 9
rect 33 6 34 9
rect 29 4 34 6
rect 36 9 43 12
rect 36 6 38 9
rect 41 6 43 9
rect 36 4 43 6
rect 45 9 52 12
rect 45 6 48 9
rect 51 6 52 9
rect 45 4 52 6
<< ndc >>
rect 9 6 12 9
rect 16 6 19 9
rect 23 6 26 9
rect 30 6 33 9
rect 38 6 41 9
rect 48 6 51 9
<< ntransistor >>
rect 13 4 15 12
rect 20 4 22 12
rect 27 4 29 12
rect 34 4 36 12
rect 43 4 45 12
<< pdiffusion >>
rect 29 24 34 25
rect 29 21 30 24
rect 33 21 34 24
rect 29 19 34 21
rect 38 24 43 25
rect 38 21 39 24
rect 42 21 43 24
rect 38 19 43 21
rect 47 24 52 25
rect 47 21 48 24
rect 51 21 52 24
rect 47 19 52 21
<< pdc >>
rect 30 21 33 24
rect 39 21 42 24
rect 48 21 51 24
<< ptransistor >>
rect 34 19 38 25
rect 43 19 47 25
<< polysilicon >>
rect 27 32 38 33
rect 16 31 22 32
rect 16 28 17 31
rect 20 28 22 31
rect 27 29 28 32
rect 31 29 34 32
rect 37 29 38 32
rect 27 28 38 29
rect 8 25 13 26
rect 8 22 9 25
rect 12 22 13 25
rect 8 19 13 22
rect 16 25 22 28
rect 34 25 38 28
rect 43 25 47 27
rect 16 22 17 25
rect 20 22 22 25
rect 16 21 22 22
rect 8 16 9 19
rect 12 18 13 19
rect 12 16 15 18
rect 8 15 15 16
rect 13 12 15 15
rect 20 12 22 21
rect 34 17 38 19
rect 43 17 47 19
rect 27 12 29 14
rect 34 12 36 17
rect 43 12 45 17
rect 13 2 15 4
rect 20 2 22 4
rect 27 -1 29 4
rect 34 2 36 4
rect 43 1 45 4
rect 16 -2 29 -1
rect 16 -5 17 -2
rect 20 -5 23 -2
rect 26 -5 29 -2
rect 42 0 53 1
rect 42 -3 43 0
rect 46 -3 49 0
rect 52 -3 53 0
rect 42 -4 53 -3
rect 16 -6 29 -5
<< pc >>
rect 17 28 20 31
rect 28 29 31 32
rect 34 29 37 32
rect 9 22 12 25
rect 17 22 20 25
rect 9 16 12 19
rect 17 -5 20 -2
rect 23 -5 26 -2
rect 43 -3 46 0
rect 49 -3 52 0
<< m1 >>
rect 17 31 20 32
rect 9 25 12 26
rect 9 19 12 22
rect 17 25 20 28
rect 17 21 20 22
rect 24 29 28 32
rect 31 29 34 32
rect 37 29 38 32
rect 24 18 27 29
rect 9 15 12 16
rect 16 15 27 18
rect 30 24 33 25
rect 9 9 12 10
rect 9 5 12 6
rect 16 9 19 15
rect 16 5 19 6
rect 23 9 26 10
rect 23 5 26 6
rect 30 9 33 21
rect 39 24 42 25
rect 39 20 42 21
rect 48 24 51 25
rect 30 0 33 6
rect 38 9 41 10
rect 38 5 41 6
rect 48 9 51 21
rect 48 5 51 6
rect 16 -5 17 -2
rect 20 -5 23 -2
rect 26 -5 27 -2
rect 30 -3 43 0
rect 46 -3 49 0
rect 52 -3 53 0
<< m2c >>
rect 9 6 12 9
rect 23 6 26 9
rect 39 21 42 24
rect 38 6 41 9
<< m2 >>
rect 38 24 52 25
rect 38 21 39 24
rect 42 21 52 24
rect 38 20 52 21
rect 8 9 42 10
rect 8 6 9 9
rect 12 6 23 9
rect 26 6 38 9
rect 41 6 42 9
rect 8 5 42 6
<< labels >>
rlabel ndiffusion 46 5 46 5 3 dt
rlabel pdiffusion 48 20 48 20 3 dt
rlabel polysilicon 44 13 44 13 3 df
rlabel polysilicon 44 18 44 18 3 df
rlabel ndiffusion 37 5 37 5 3 GND
rlabel pdiffusion 39 20 39 20 3 Vdd
rlabel polysilicon 35 13 35 13 3 dt
rlabel polysilicon 35 18 35 18 3 dt
rlabel ndiffusion 30 5 30 5 3 df
rlabel pdiffusion 30 20 30 20 3 df
rlabel polysilicon 28 13 28 13 3 wt
rlabel ndiffusion 23 5 23 5 3 GND
rlabel polysilicon 21 13 21 13 3 wf
rlabel ndiffusion 16 5 16 5 3 dt
rlabel polysilicon 14 13 14 13 3 Reset
rlabel ndiffusion 9 5 9 5 3 GND
flabel m2 38 20 52 25 0 FreeSans 11 0 0 0 Vdd
flabel m2 8 5 42 10 0 FreeSans 11 0 0 0 GND
flabel m1 9 15 12 26 0 FreeSans 11 0 0 0 Reset
port 3 nsew
flabel m1 17 21 20 32 0 FreeSans 11 0 0 0 wf
port 4 nsew
flabel m1 16 -5 27 -2 0 FreeSans 11 0 0 0 wt
port 5 nsew
flabel m1 24 29 38 32 0 FreeSans 11 0 0 0 dt
port 6 nsew
flabel m1 30 -3 53 0 0 FreeSans 11 0 0 0 df
port 7 nsew
<< end >>
