magic
tech sky130l
timestamp 1636602913
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 10 20 12
rect 15 7 16 10
rect 19 7 20 10
rect 15 6 20 7
rect 22 10 27 12
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
rect 29 10 34 12
rect 29 7 30 10
rect 33 7 34 10
rect 29 6 34 7
<< ndc >>
rect 9 7 12 10
rect 16 7 19 10
rect 23 7 26 10
rect 30 7 33 10
<< ntransistor >>
rect 13 6 15 12
rect 20 6 22 12
rect 27 6 29 12
<< pdiffusion >>
rect 8 23 13 34
rect 8 20 9 23
rect 12 20 13 23
rect 8 19 13 20
rect 15 19 20 34
rect 22 27 26 34
rect 22 26 27 27
rect 22 23 23 26
rect 26 23 27 26
rect 22 19 27 23
rect 29 23 34 27
rect 29 20 30 23
rect 33 20 34 23
rect 29 19 34 20
<< pdc >>
rect 9 20 12 23
rect 23 23 26 26
rect 30 20 33 23
<< ptransistor >>
rect 13 19 15 34
rect 20 19 22 34
rect 27 19 29 27
<< polysilicon >>
rect 20 45 25 46
rect 20 42 21 45
rect 24 42 25 45
rect 11 41 16 42
rect 11 38 12 41
rect 15 38 16 41
rect 11 37 16 38
rect 20 41 25 42
rect 13 34 15 37
rect 20 34 22 41
rect 29 39 34 40
rect 29 37 30 39
rect 27 36 30 37
rect 33 36 34 39
rect 27 35 34 36
rect 27 27 29 35
rect 13 12 15 19
rect 20 12 22 19
rect 27 12 29 19
rect 13 -4 15 6
rect 20 -4 22 6
rect 27 -4 29 6
<< pc >>
rect 21 42 24 45
rect 12 38 15 41
rect 30 36 33 39
<< m1 >>
rect 12 41 15 51
rect 21 45 24 51
rect 21 41 24 42
rect 12 37 15 38
rect 30 39 33 40
rect 30 34 33 36
rect 9 23 12 31
rect 22 23 23 26
rect 26 23 27 26
rect 9 17 12 20
rect 24 22 27 23
rect 30 23 33 24
rect 15 11 18 14
rect 30 15 33 20
rect 39 17 42 51
rect 9 10 12 11
rect 9 5 12 7
rect 15 10 19 11
rect 30 10 33 12
rect 15 7 16 10
rect 22 7 23 10
rect 26 7 27 10
rect 15 6 19 7
rect 24 5 27 7
rect 30 6 33 7
<< m2c >>
rect 9 31 12 34
rect 30 31 33 34
rect 24 19 27 22
rect 9 14 12 17
rect 15 14 18 17
rect 30 12 33 15
rect 39 14 42 17
rect 9 2 12 5
rect 24 2 27 5
<< m2 >>
rect 8 34 13 35
rect 8 31 9 34
rect 12 32 13 34
rect 29 34 34 35
rect 29 32 30 34
rect 12 31 30 32
rect 33 31 34 34
rect 8 30 34 31
rect 23 22 28 23
rect -12 20 24 22
rect 23 19 24 20
rect 27 20 48 22
rect 27 19 28 20
rect 23 18 28 19
rect 8 17 19 18
rect 8 14 9 17
rect 12 14 15 17
rect 18 14 19 17
rect 38 17 43 18
rect 38 16 39 17
rect 8 13 19 14
rect 29 15 39 16
rect 29 12 30 15
rect 33 14 39 15
rect 42 14 43 17
rect 33 12 34 14
rect 38 13 43 14
rect 29 11 34 12
rect 8 5 13 6
rect 8 4 9 5
rect 0 2 9 4
rect 12 4 13 5
rect 23 5 28 6
rect 23 4 24 5
rect 12 2 24 4
rect 27 4 28 5
rect 27 2 48 4
rect 8 1 13 2
rect 23 1 28 2
<< labels >>
rlabel ndiffusion 30 7 30 7 3 Y
rlabel polysilicon 28 13 28 13 3 _Y
rlabel polysilicon 28 18 28 18 3 _Y
rlabel ndiffusion 23 7 23 7 3 GND
rlabel pdiffusion 23 20 23 20 3 Vdd
rlabel polysilicon 21 13 21 13 3 A
rlabel polysilicon 21 18 21 18 3 A
rlabel ndiffusion 16 7 16 7 3 _Y
rlabel polysilicon 14 13 14 13 3 B
rlabel polysilicon 14 18 14 18 3 B
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 20 9 20 3 _Y
rlabel pdiffusion 30 20 30 20 3 Y
rlabel m2 33 2 36 4 8 GND
rlabel m2 36 20 39 22 7 Vdd
rlabel m2 36 2 39 4 7 GND
rlabel m1 21 46 24 48 5 A
rlabel m1 12 46 15 48 4 B
rlabel m2 39 14 42 16 7 Y
rlabel m1 39 46 42 48 5 Y
<< end >>
