magic
tech sky130l
timestamp 1636167701
<< ndiffusion >>
rect 8 13 13 16
rect 8 10 9 13
rect 12 10 13 13
rect 8 6 13 10
rect 15 6 20 16
rect 22 14 29 16
rect 22 11 24 14
rect 27 11 29 14
rect 22 10 29 11
rect 33 15 38 16
rect 33 12 34 15
rect 37 12 38 15
rect 33 10 38 12
rect 44 15 49 16
rect 44 12 45 15
rect 48 12 49 15
rect 44 10 49 12
rect 51 10 54 16
rect 82 15 87 16
rect 82 12 83 15
rect 86 12 87 15
rect 82 10 87 12
rect 22 6 26 10
<< ndc >>
rect 9 10 12 13
rect 24 11 27 14
rect 34 12 37 15
rect 45 12 48 15
rect 83 12 86 15
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
rect 29 10 33 16
rect 49 10 51 16
rect 54 10 82 16
<< pdiffusion >>
rect 25 29 29 33
rect 15 28 20 29
rect 15 25 16 28
rect 19 25 20 28
rect 15 23 20 25
rect 22 28 29 29
rect 22 25 24 28
rect 27 25 29 28
rect 22 23 29 25
rect 33 28 38 33
rect 33 25 34 28
rect 37 25 38 28
rect 33 23 38 25
rect 44 27 49 29
rect 44 24 45 27
rect 48 24 49 27
rect 44 23 49 24
rect 51 23 54 29
rect 68 28 73 29
rect 68 25 69 28
rect 72 25 73 28
rect 68 23 73 25
<< pdc >>
rect 16 25 19 28
rect 24 25 27 28
rect 34 25 37 28
rect 45 24 48 27
rect 69 25 72 28
<< ptransistor >>
rect 20 23 22 29
rect 29 23 33 33
rect 49 23 51 29
rect 54 23 68 29
<< polysilicon >>
rect 63 51 70 52
rect 63 48 66 51
rect 69 48 70 51
rect 63 46 70 48
rect 15 40 22 42
rect 15 36 16 40
rect 20 36 22 40
rect 15 34 22 36
rect 44 38 49 39
rect 44 35 45 38
rect 48 36 49 38
rect 48 35 51 36
rect 20 29 22 34
rect 29 33 33 35
rect 44 34 51 35
rect 49 29 51 34
rect 63 31 66 46
rect 54 29 68 31
rect 78 27 84 28
rect 78 24 79 27
rect 82 24 84 27
rect 13 16 15 18
rect 20 16 22 23
rect 29 16 33 23
rect 49 16 51 23
rect 54 21 68 23
rect 78 22 84 24
rect 78 18 81 22
rect 54 16 82 18
rect 29 6 33 10
rect 49 8 51 10
rect 54 8 82 10
rect 13 -6 15 6
rect 20 4 22 6
rect 29 5 36 6
rect 29 1 31 5
rect 35 1 36 5
rect 29 0 36 1
rect 8 -7 15 -6
rect 8 -10 9 -7
rect 12 -10 15 -7
rect 8 -11 14 -10
<< pc >>
rect 66 48 69 51
rect 16 36 20 40
rect 45 35 48 38
rect 79 24 82 27
rect 31 1 35 5
rect 9 -10 12 -7
<< m1 >>
rect 65 51 81 52
rect 65 48 66 51
rect 69 48 81 51
rect 6 36 16 40
rect 20 36 21 40
rect 78 40 81 48
rect 24 28 27 39
rect 45 38 48 39
rect 36 28 39 32
rect 45 34 48 35
rect 69 28 72 37
rect 78 36 90 40
rect 9 25 16 28
rect 19 25 20 28
rect 9 24 20 25
rect 24 24 27 25
rect 33 25 34 28
rect 37 25 39 28
rect 33 24 39 25
rect 9 13 12 24
rect 36 16 39 24
rect 33 15 39 16
rect 9 8 12 10
rect 6 4 12 8
rect 6 1 7 4
rect 10 1 12 4
rect 6 0 12 1
rect 24 14 27 15
rect 33 12 34 15
rect 37 12 39 15
rect 45 27 48 28
rect 45 15 48 24
rect 72 27 83 28
rect 72 25 79 27
rect 69 24 79 25
rect 82 24 83 27
rect 69 23 72 24
rect 87 16 90 36
rect 0 -7 13 -6
rect 0 -10 9 -7
rect 12 -10 13 -7
rect 24 -10 27 11
rect 45 5 48 12
rect 81 15 90 16
rect 81 12 83 15
rect 86 12 90 15
rect 81 10 90 12
rect 30 1 31 5
rect 35 2 48 5
rect 35 1 51 2
rect 42 -2 45 1
rect 48 -2 51 1
rect 45 -4 51 -2
rect 84 -8 87 10
rect 81 -10 90 -8
rect 21 -11 84 -10
rect 21 -14 24 -11
rect 27 -13 84 -11
rect 87 -13 90 -10
rect 27 -14 90 -13
rect 21 -16 30 -14
<< m2c >>
rect 24 39 27 42
rect 36 32 39 35
rect 45 31 48 34
rect 69 37 72 40
rect 7 1 10 4
rect 45 -2 48 1
rect 24 -14 27 -11
rect 84 -13 87 -10
<< m2 >>
rect 23 42 28 43
rect 23 39 24 42
rect 27 40 28 42
rect 68 40 73 41
rect 27 39 69 40
rect 23 38 69 39
rect 68 37 69 38
rect 72 37 73 40
rect 68 36 73 37
rect 35 35 40 36
rect 35 32 36 35
rect 39 34 40 35
rect 44 34 49 35
rect 39 32 45 34
rect 35 31 40 32
rect 44 31 45 32
rect 48 31 49 34
rect 44 30 49 31
rect 6 4 12 5
rect 6 1 7 4
rect 10 2 12 4
rect 10 1 21 2
rect 6 -2 21 1
rect 42 1 51 2
rect 42 -2 45 1
rect 48 -2 51 1
rect 18 -4 51 -2
rect 18 -6 42 -4
rect 81 -10 90 -8
rect 21 -11 84 -10
rect 21 -14 24 -11
rect 27 -13 84 -11
rect 87 -13 90 -10
rect 27 -14 90 -13
rect 21 -16 30 -14
<< labels >>
rlabel ndiffusion 34 11 34 11 3 #6
rlabel pdiffusion 34 24 34 24 3 #6
rlabel polysilicon 30 17 30 17 3 out
rlabel polysilicon 30 22 30 22 3 out
rlabel ndiffusion 23 7 23 7 3 GND
rlabel pdiffusion 23 24 23 24 3 Vdd
rlabel polysilicon 21 17 21 17 3 in(0)
rlabel polysilicon 21 22 21 22 3 in(0)
rlabel pdiffusion 16 24 16 24 3 out
rlabel polysilicon 14 17 14 17 3 in(1)
rlabel ndiffusion 9 7 9 7 3 out
rlabel ndiffusion 83 11 83 11 3 GND
rlabel pdiffusion 69 24 69 24 3 Vdd
rlabel polysilicon 55 17 55 17 3 Vdd
rlabel polysilicon 55 22 55 22 3 GND
rlabel polysilicon 50 17 50 17 3 #6
rlabel polysilicon 50 22 50 22 3 #6
rlabel ndiffusion 45 11 45 11 3 out
rlabel pdiffusion 45 24 45 24 3 out
rlabel m1 81 37 81 37 3 GND
port 16 e
rlabel m1 9 5 9 5 3 out
port 19 e
rlabel m1 9 37 9 37 3 in(0)
port 20 e
rlabel m1 0 -10 3 -6 3 in(1)
rlabel m2 54 38 57 40 1 Vdd
<< end >>
